��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� rā�SZ )����C.��&0C]�-��[�3�-���+��պݣ�k�J�vo`�A�����f����u�X���v�=�а���]Q�Wۿ�߸�=_Q�X����j>��Zw�K��SvX��ƥ.���#�����Z�0���#7{��\S$��@1I�QX~TQ�E��db����۰� ���>0�%�9�j汈��}��1� ��2���h�G��SeY�a���	'<x�p��k�H`�H�j^y�0�s�78+���ֳ�`�R3dW��_��{p[�?$�s0��#�zS�_��bH
�c�p�IL7]� |����Q�� ��Rr���=��E즕2%�����`�^��l�q-�]�p��jf��Ӽ-f%H���ȳ�>��+���M�71��4_�) 3�46h�rb�J�W� k�h~K0�>P$�_n)���5�r�j��W�J&޴o��$>��6��ŀ�;A~<6P��K�~��f��*I
�Z��}`q���ApC��n���g���3��-�іrO�mF���,�$��@�BI�q�}��Ȥ֐����î�䂧��@������U���vU������ �T#K@f�㯁����|95<@���+�-�)�����K���FI�k���*@�m&���
���ma1[�2�u�I�\�U�yu���o�|��2����;�W�W�}P�K>%5�'�8���׫=����k��,�t�M�0�8]q3���N���GvZ�A����^�Љ'r�n�yG�pI3Vu�ҶU
=��� �Ï·lqo�P�!����P�����^pHw]��*�
�~�w��l�.#��D��fZd�6���zd�M������R3v"\�������4Ӛ4Θ��lu�A�ٓ�';�w�X��XD���{����7ƔIWrK��
�*�/��J�׍d$�����r�ҹbWA6U�U��Ŏ��,��<�3	��l{�ځaϚ��~Tt#����|�������}n����<�+�oV�&?�e�{�q~�Sz�l$��}TQ�9!Q�_f�kH�,���B�#C*���Xjƿ�]�)�k�Z�=B �
a=���S�#����.�}=$�.�Cc��(�����<�x������2�z��E=�v=���S�y�Jf�}��wĖ+��	�O�Ps����פP#�i��9+��l���/u�W	��\�[��.������}9�Z�R$ym��y�ׄ*W�D��%�\�҉*�!(�9Ҹ&/��o6%ԃ��= WZt����?V��Q&�j��U��~r[�����JB9t`�QSH>�7S�=�E��h"٢c���M�;��	]Pil!$I�e#�K�Gs�x�U�Pprfy��Y�\j�2��69��1*!��ll��~�}$NEғ����O�^t>��dk9���?�\8�Y��Q͑�"���X3��f��'�~�jR��ױ?T^qT�wN3e�TZ�(؄�>�������ߐr�0�]C��s%Y	�-����#��
���UVnV:@g��H8ޔC��f��u��!Fƙstʫ_t��� ��߳xQ�-)�\���#��Fv�d x<��iA�v���u�#�"�I6s��H�q��D��l� �J��*�(��^շȅo��ywγ@���n%�(�m$��j L�kHJ�/��`S�R��U�������g*0`?��%��xQ\��� �t-��6܃���~S�vϡ�&��R[�)��5u�WnG۬����R��қ� �@[I|N)q���[�n��Y���)˅xJDȕ֫e�*�>��$�������q�����o�1���4$���N�cɞ�x������L��d���j�����r�@W����Mxi�F�M�7��LB�U���=�'��-�6�����{_!����G<�"ҹ»���~��/���jA�M�JH�E���[��&���A��HxW��� ��X5�ힵc#b�|)����x�(�rxY��Ѧ�m^m�l�C��t��=*ל�Xy9�r�YN/��G�����!=���p	��%�O��e��Z,��zu����"��BM���]b��!�T��N�ru�����:�nz<�>��b>��\�z�T�)��Т�W ��N�b�P%8����w�*���@���!��ue�J��}�C�f�^I̥��_�[K"w��\	�O�Z���?y�x�K>��(j��M�ӉH�C	+�%�`�)JM�o9 h��g�Z0ר��pN�{]8�6dBN�&��f����;R��������mڿ�^�}-4�jѳX>čEv�*����zf����oT���ЬC�K��v,K�g�$3��֯j�k��Tt���/߂I��X����Yo���BEZ���!V1�3b�9���C�i��BȄ�Ʒ��=�'�%�����d`-%I�RJ P�������r�⢦k�\6"��ئ}���Ο����+-˪���F�5?%���P��f)Xj�j��!BXJԊ��#φ�^j���}��P([9���d$<{� �׿$�5e����J��Y'CVh���H��3��V?���%,W8����{H 1t۞�l�]��ɠ{�_�w���Z�e���8��#�6�6�q��&���df�=�y�ì�C��[�ͧ����������\M[�U�B<� �/����uh���OLVr��_���#Q��p��!�#PV����l�
'�CƵ�K�z��b�s�Z?���-��<�'�2J �����'���z�e'�n�%J��2�a�4�T(��7?���bU2��l�?��o^�Y���I	�_������Z�s$�%M�(�#Ǎ�m��}$m�� 5Qk��fft37nM ����5l�ᨗ����MH�T=��1x*�l��_V�ܾ=��m��u�8G����I�J+������ ���0&p����俠��|�UA=�\ʐ^�P�I��}K��E�t�B�*��a[�����[.ۡ�ڙLM;�,���t0��\$R�8�]�ּu�F*����0,ӂ=���mR}u��t�H𙑏#}5��v��T-�n��K\0S���Ϣ����ٍ�I�%��U�f�t0��&J2�s�L=ֺZT�	
�E��)�[�+�{ø4$2J�ꊥ�7����\f��;d��C@`.l��>Xz�!k�c�d��ȕk����E��C�p��(,����GY��+�Ƚ?[�Ƙ=����Gu��!�==�U�>� �!?�:(_�3�@kÒ��E�x���Z8��P����L[��'��Tކ�0k��l��@|�y�c�M"�h���" }������R*]�Dn����I
?%@�����Y�"�8a)���ʄ26E�;�'[(�`lh�b|ҕ���2�����|�#"