��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� rā�SZ )����C.��&0C]�-��[�3�-���+��պݣ�k�J�vo`�A�����f����u�X���v�=�а���]Q�Wۿ�߸�=_Q�X����j>��Zw�K��SvX��ƥ.���#�����Z�0���#7{��\S$��@1I�QX~TQ�E��db����۰� ���>0�%�9�j汈��}��1� ��2���h�G��SeY�a���	'<x�p��k�H`�H�j^y�0�s�78+���ֳ�`�R3dW��_��{p[�?$�s0��#�zS�_��bH
�c�p�IL7]� |����Q�� ��Rr���=��E즕2%�����`�^��l�q-�]�p��jf��Ӽ-f%H���ȳ�>��+���M�71��4_�) 3�46h�rb�J�W� k�h~K0�>P$�_n)���5�r�j��W�J&޴o��$>��6��ŀ�;A~<6P��K�~��f��*I
�Z��}`q���ApC��n���g���3��-�іrO�mF���,�$��@�BI�q�}��Ȥ֐����î�䂧��@������U���vU������ �T#K@f�㯁����|95<@���+�-�)�����K���FI�k���*@�m&���
���ma1[�2�u�I�\�U�yu���o�|��2����;�W�W�}P�K>%5�'�8���׫=����k��,�t�M�0�8]q3���N���GvZ�#z�HM���f5�����;�q��Pj����H�L�}��T7���z@�o	%�PFmy�lc�
)�8yIf�o���Z�"4��r���o�6˦��)��"�~���6��}�pY���]��
��K,�	���1D�̹�@��$���(_kk<| &���x,�u��Sm��Fģ	U��U9�k-��c�KU ��1$k�):h�����!�Έ>�l�B2A�V쉀�#� o�Aڐu�Q�%`��ܸ��cb.�����E��&�Ѯbz-V*�E���bnjۜb>W���z�<\UlA"���i��J��Xj݊���	p��k��1O:�$w%�C�\��H��U���Z�W��k�B�E��d��/���|�0�=o�g����/Z^����X@�N �Y*E�M��j��Ʒ�G��V��$��Qhw-J���,�B�����>�n�N9+���̍�)ТP��yw�~2�]�4�E�,��$&�_�������%�#P� M����PA��[�Z]�ϒ=!�ܠ��T�X�`2s��gq�D���&��%�?�Gy���4E��[4�͹��*�r�S�Q�����!P<�g����j�m2W|���i�:�?���_7��[�@k��v��I�������,��u�T�䷏Cë(��5<-�����8J���R�[{{l�Ijt�d�	0�:�K���}�� ��@W���D���&�b�kݿQ<
�d�dl�\aJ�n��En�V���pT���u!=��$�Z�
���Ѭ�!���w�*� ���NثE�_ *X��F�A
^�7��u ��*r�ܜK	���7�,+�iպ��z��<�7��x�j�ԡ��ܿ�bx2w-�lvDd�T���$:�k��l��Mr �n诗�Tcpb������/��h&�=��|�B"����Yb�=���t-�B��[K߹�zKVX�ʳ���_N��hF�Z�3 �<�~[0��s�ـ�`��=B�:��p�C��O#`z�&7a�Ђ����Z�2 ��=���Ṉ���ҙ�ѧ���q1��E�nMS��E��n�E�&�V���Y!S�ҍLIW��:��Sǥӱ `�,a!H����F�W��_�54������dPu-���
LU�ܧ�ljy�}���`̒�{+�W3<��N�//~�d���M��v�f�a����"���OA��>�#���t���������Z!QL�'�@�"�g��������W|���+Xfg*�Рr��u/��B96IWX��t�з���l�.����p�u�S���T��@p�v�m�2���m�#3�]G/n����BJ')0����
HD��� �[_+��u؁)�t����r��٤�}�2ٿ����+Qj�����S���|b�$�F];����U��",!��&�$��`�m��<��n����'E�\�����_kջRh��)��I�х#n�{�����[6d��/YhW�*Ѡ�iǏ%zB�
�U]~-|��U���ȩ�i���hD�ZӞ�sM�a6�f�4Ľ��`|�W��(��B��7ppHO&�:�P�I�r�<��t��S��n5˟��ˇN��p|��#~1'�J��E�{��$�5�������]�Y�^��r ���?�WH��w5f�˒��;�H܊Y-8FLn�������|ۻ�"�K��W ~� :l��D��tD�B�%��A���̅�
��.�(�t����,�C���A��4�=Q�`8bQ�whE��k�t�]�"�G��A�����*��J��*�����q����9Ec�Yi%X�a4�;�Sn�R҄�`�Lf�ɨ�Ԛ	�G	Y{0혗T5�p7�F��<Ès��ȕ	����������%ᢨ��!�Do2��m�[g�����\�������G��h=;}���m���Ae��GS+s��F��l*�p�ʘ���J����M�v �xB�����+�ʲ)N��H|=�5&0]ގ'gP����>�����EW#��w�n�y��aی�2��3tYb�ƻf��?P>��*��Z��~���wI�ߕ,Ӱ�*���0�M%��O�J+��&��0�;
}}#K�i���(3t��ÅHW)�k̫ �/<���ӧ����K��u����)���^���3J�)�@���J��Pu3�\A'��, �R��h΅�*n�����5�l� ��کn�u @o�F7��.�2=���[�7��$��`�$F����S�#4�� sN��G^�5�	q�]�1Jx+��U�m�6p���|~�Nآ�Z�?�{L�2'<��uc؀n�a��������WGz:��܎c\MA�5@|�Tc��a�	���uv�L
�uS�%.��k.p[*�ֵ�	wu}�,6���>� �542��Ql5�� �y���j:'������Y~�!��.,��r3Q�.��/�>f���!��!�ȷ�b�H�qtG2��U�N�w��A���\#�r�U�\�)R�\!�N��UT
���tŰ�k@�El�,�@�9P}L�]�6�r3ʿ����wTŎ�;/����_���+3��Zu�R�Qߪ�Ȫא���W�Om��Gu�	-w�hO��em�q����~@�h۶8��wk�BU��a�ß���������>�-J��îf2}y�����"��ｏ�Ig��S�/v��%��L�%w������Q�E<q�/��}c�\�x�P�Jj+Aw��SHѴ������N�Bɮ%�}���p'�fa����`�_�AZNj7卮������ W6ٿ�~f.��9��Y�/w<G�9���mC���#Z:~\� jə-J�ǜci��<�p�U}2�Պ9Z��4b�jB�������k 1��-g���5�7��]���k+p��&��e�]�����P����a��o�P��7:�s��o�5�H٣Z�XS���%hx��R�ت�̈,��#�4��,_�(0ANB��YŵB�<�&�KDɿ\~@��'�w&[>)Ì���#���I/T�0�"g���x�]�?���
�
�#� [��_����fn
x��"C�p�l�9�,�,��cF�v���y���W2�^�O�mQhTϞv'����Db��r�_�!�#}�aٜW��o4/�,^ll�U���^�}άmYv�p۬�F�lO�� �l�m�l1EM�I�a�{�l�C;^ø�	�26,�灛����<��J�HC��Q���b>x�m� @8)
��)u�B�,q)GJ��VU�d$|h<|4��) �+��T��c歊�A��4q�6t��l�#�ꗅ���)@[\���L�{o��Ǟ���&�K¡`�o��I��[����w#z%�*�?s�0�1ek�� ǲ��>g�z���;���K3'D_4��X�	�q�8��J�Λ�EǷ3��k z9P����8h1[��1� ��9^4e��� g^X;�\��D0�߸wU�1Ck���	,�#�0&� G�ww�\�>����{�n�!��}G�/L��Z����(����q��=��A���U�,�	L��*���z���D�L�A�s~0���ԸK��P�"隮��%Q�K\�w� ׾?��������Csj��t����0*џ����͹�e:6�A�VduG%���#3�?�#َ�������/�S���ɰN^M�AyZ) *
��fu��_��/�}Y���������95M��$�il;�L.����b��~���nq|��W��+�f��<�Z�]$����>jTԬ�����W����}�X�+���=¾���(�Q��F�B�����؅yE�����2��tCA(n��]�/V�̈
�G��Z�Č �h$�.6qo��_ޔ�^6070.��t	�XB�G��N~��N,���V{�: ��!�VrR>��;�ѐ��qk��2�}r���l�MB�̳��bi��n* � �ʾ�L��_�˼CE��~�t7�@��J�Mft����\�b��~���l.���h��Z���,��6�z#&`\xN8D�^t~�ZϹ�|�wZ$���M��C��e3�z[�Aq(X5h4���V[���̏�;5��1|[;%�i%�m� ��Z&>ԋ���u|H�֬��Ʈ�r�w&.c!A)X�6V$<~��N���L2T��wO����J���|˧�$����Z���鞜����ϊ�q�dg�:%t��D�3\IsW�\�v����?�*��������a�u|�N=Y)h�����V_)���ڗ����O�I^���d����j� �J5�$"ވ������t�r7�VŕH���\2�٣����H��4w�V8�A׹aU�-�.�Z�����R���3�	�{�VhÈ�|�k��WѾ�"��ɏ�z��Bѵ�_&�����p�a탷���V�I\6R��' P)���2�B�� ��"!欏�dD&%��<K${��,F���6��!����'�:�=w1�_n`'?�+�&�d.��L:��k)��Է��
�˓��/��9�\��/kr�F� TM��MY�Ns}��+�@\�Qx��,˘��6��H�o��3�k�;dց�`�T5{m2�CVocй�/����E9J�:d��'W���5�����V!=��9W۠΀������qRMʗɞ�BrT�~�,��M>�v_�v닔2��Z;b8�A0G�'�} o;�0~��Dw����&}��gs�z�U��2b��l
8���1�wHC薁Y[��