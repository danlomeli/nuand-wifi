��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� rā�SZ )����C.��&0C]�-��[�3�-���+��պݣ�k�J�vo`�A�����f����u�X���v�=�а���]Q�Wۿ�߸�=_Q�X����j>��Zw�K��SvX��ƥ.���#�����Z�0���#7{��\S$��@1I�QX~TQ�E��db����۰� ���>0�%�9�j汈��}��1� ��2���h�G��SeY�a���	'<x�p��k�H`�H�j^y�0�s�78+���ֳ�`�R3dW��_��{p[�?$�s0��#�zS�_��bH
�c�p�IL7]� |����Q�� ��Rr���=��E즕2%�����`�^��l�q-�]�p��jf��Ӽ-f%H���ȳ�>��+���M�71��4_�) 3�46h�rb�J�W� k�h~K0�>P$�_n)���5�r�j��W�J&޴o��$>��6��ŀ�;A~<6P��K�~��f��*I
�Z��}`q���ApC��n���g���3��-�іrO�mF���,�$��@�BI�q�}��Ȥ֐����î�䂧��@������U���vU������ �T#K@f�㯁����|95<@���+�-�)�����K���FI�k���*@�m&���
���ma1[�2�u�I�\�U�yu���o�|��2����;�W�W�}P�K>%5�'�8���׫=����k��,�t�M�0�8]q3���N���GvZ�i�+ C�e
��Ќ�S�v<%���q��e_��
�k�夞��>ZO7E~��5k�TW Aod��eE���G���ɑ-'���?�G$����ќ����8ɸ+ 5ʗ���l�d��,�J�
�^�3b,�����J����#n�zK����z�&��;|�\�^���'e�W�����">�w*	FO�Δ��v���I�h������l[�tgOy \��\�<�ʏz�V��<CwR0NgE1�.�����!�]�q�'P�B��!��		?������_��'��_Xh��<�*��'�BJeg�+@囐"��Bz��
~&e�ͥ��߄|�X9���-�7G$�	��V((�d�e���5
E��5���pz	����v �z[����$�^՟��s)X���F�P���0mv�귲��b4]�'[�d]�.��FW�n�(��&o�*Յ7��})��O�]7y����C��z9g��pr���wD�p��y`I|����t��@OSz��w	�K����7��ӁC@���`hK��=g��I?SR=�+dx9]��t��,(	u4rƇs�|��C��|��u��}��b�Pz-�����cB���������3�6�	��F��H��w#��C�j�,��	)�(�DF�P�YB̐��-6��J�my�>�������d�������'����㸽��;��	E8#�{�l�h�,�Ȧ�q�p�8��?t��n�G��ylB��Al��c�z.��x�s�yG�A��G�H/�L�2(�Uf|z.�\������JR&�/�j�;1�`��\���m;^ �����:�O��n<�� }fm�	��ڏ��^��H�A�t�e��Y"U5��ު;'}<�����TzV��Ո�����o'����}1�w�QJϧ*�F�.`����&z��#��E+��Ƭ���$ �3 P&XJ�:����ׯz����2���U#l
�lJ�dW�n���Ϋ�G�\�����zw=��C?����y�9��Z�XYp��F�py�U���W��K�]�4�������9�G�޽���p��h,*Lq�~qi���!u���'�j$�ayEs#/|�Z�`V��󓘱�5Y�����z�!`c߷x�b���$Y5?V>�ˇ�.�I�"�'JZx���
g��F�J n��S�*�����؍�k�0�M5L������4X�����C���u�$7@�֥ʅZ-��R��	�V,�)�8}�7�(fM�m�$�ety�⾗���AH����`�G���J���t&Ѱ���巟��*zc�_���K!�e5<��ï����D������0+z� �m��6�S���y��[����*��*(|@���?m\���b���Q0�wW�0 3X2��������ꜷ3���VTI}eͦ\�v��Aw-#d����������9_��.p���7�+�>�xT*��30�Y�M�<��
Ţ"�a�mJƷ7�6���Alim��946%�c6�Zs&�_�H��7��>ɧ5v��=��5ۉ�%.x׎^Eq�YE)����8,�t��K���uPk�;ˠǮ|X:De��P��0q�C��˳�a��Ԓ���ӛ!�*ʯ:��5�����Šj�+��z�ǁ$�<�ȣz�`��8�OYB��IM��D h��7e����=Q�5�k����,E� ��Ѓ��$1͈b�ޒe���MwK��,�p��W�M�|%���7��!z�)\T���	�EU@�T�7x�#����Fc��F�>�+g�q�8��-���� �~��A��c��D�,X�=���|�!�ucZ���ѹ�N+{�=�@5Gd�����!"~qΤ"�D�d|����<����~�x-�|��`C�
�|�ֺx��X��r!�~�����KL�1�� WXF>�ٞ��r���Py
�H�D�?�{���c�E�j5�R�LK�\&&�Bfm@��**�ܩ̆[0,�o��YzAk�y�a(#�*j�VN���)b��c��i}7o��]ϧM�D�3z*��?��~x�E�M�E��'�����lqiw����!��1ѱ�zJ�^��� w��~���3I%�����;p����we@UXhoMf�mz�Y~��z�H����+\��
\p	C�5B��g��?R5�Y�Hس���qC��k�{E«Xb��$�$�B�}�)P��**ړ;>�]v<7Ҡq�O�/E9�l&�J�;�� �Ol�9�B�2;��i����еx��|x�0(�O���ߴ�*5D���"��-;�R����|�P������/Mmu }��@m���K���8o�q��A�sR2��A;.e����2�6��!�tYwT�x�'���?�N�����\�S�5��l�@8�[hCoݫ̮c$
S�ĠA����c��͵>�Y����l]ͻ�=��\��b��Z�����n,j
�o��G|w���D����{ D0��x�\�T��Gt���!��x���h����༮���@)0�u��u4d�A=�>�a��J��5�
OF���Ir�ί�(�.u,�+��#p�)����*�vΒ�5�)J��h��Cnά��N�癑��=S�C������n��*6v��l�پ������z���Q�9�:,s�I9U�뽋5���ڋ�e]��Y����KP� ?Uܙ_�[� �j����%A�H._����t�1&'+��zm1j�󼵳+h-�^6]�:Ս�L��|C��uh+lQ �W~�����hQS1z�oPaN5�4?`t%.���������F��3*��3����K$��m��e�uu��>����=��6\������'��6���Ä���5I�p���Cm9��m7�ļʺ�`��O�a���dh	M�IO��t���#��Kħ^@�*=Q��.'ۺ)G6��`l����:�s��.�B���"Gz#�OͶ��@ޓ����z��R�%vMLV��/$��Z�.�����(�D0k=[�ZG�l�j��0�,$]��35^$�n�`��^^�3��H^��<X�����W��"!�6���C���p�z�ʻ5��8]���%qelJ�`����T�A�b0ӌ�n����Gi8,6���ԛq�%�s����K�-�\�@�ՅA�a[q�l�,g�`����>L��wr�{2~�q�N��u�7��y�"n�(�&��;9���/'���c@�a�T����K8cO��
#쯇Q�:7�i;�����`���0l7���j������`/t~���X � ����p�l��t��H�˗q�F\�NQ���cد�^��_iȡ��aȻjĂ�yO��ٗ	Ǟ�:?��O��j�B)G��Z����R��0�N8C�7On�	@��?��8k�r��oJ�C^ߗ�Up�y9M}__?�_wEC3-uձ�9����|��m�T<��J�ם�����A����i��|��%�ZN������_�]J��"����WpM �<^�LK2���6�x�/[������)�r��y��|��i����y����N��goy�-��
��r����&�i���Ǧ�	����tQ(�����zLH�a�ܕA/��*�:���Ќ}��P:{�#%�l��T���B�J��$d�J��{A�(�k:��㩼�f;�_�i:߃�l���X���bX��	[���2�D`��^#�B�!���x�Yj3Z����f2	�V�0`a��Ёy2g���U�?Wia+�m6�pt>a��Y���XS:<�Zc;����d�99��F�NVs�m&}��������Ӥe�_�:&8�?�!I\8b|�7���h��������V�-��E�7N�+L,�n�����-`��V�����~p3Z|��UMր�<�&8ൺ�����1y�z/� ᮘ���(��� V䚇s��Z����3����Z����X՞4j�bU�1):}OQ4<6��Y0��E-O��Hg�`����,��\>᥉�� _$	�ѯ+4橄p�´_0�j#�o���F�{���YrsH~�P&�N�F�{MD˒I0;�ӧ|H�*�b��S�i�$4��{�8��Oti}����+u%۲%5�_#N���,{��ȷ)��6����vSѹL�^=`8ĆC�����JӉ�3�8x�����3��!RO?��� ��R�nU�[,�	�oKC$���Y\��q����ݘꬠ���(k���*`q���q�ֱ�h$$�ƪ� �����k%� GnJ�$!�ת��
��Ɩu�K�w���	r
k��χ�T�0�Wm?[�Z �����cO�'��l|l�H+EzfI���&�T���a��$��3�m�>������G���R�3i�Wȗ�e�̅`�e��M��z���>z>�/�aU��m:��S�#�	�J�_�?�������ա?}?h x��fRp�ߑ�Z�)?��c��H*�׳�^��3�k��9�j�1��h��B�G�p������2-��[��1+D�2/�>	�ec�voL �>]d�p��ոdcި�^\��U���v9�X9��(���	f*;B������8��86>��x,�=���)�,R~	�_?+�ɶ�u'Q׊���zs�L�r�UW��Q��ˊ�`{^�&��.���]c�`�u_|�%���kۘ�Z_2��"���WP���oQ���>7H `ud�Z�����&�6IԇH=�w��C�C/���K��M�7�q��d������C���Z��>?�'z�:�Z��0�7:xٚ�t`�H#��=��w�����qG�q�S�q�`Vu��q�"���7s530�v�zdu�\�G�>"�]�n����m'k�c�fF�޼�`p����oz*Yd۴�����@Q>ם��Rp��TZ;,�OaO0ۮ��V��?��3>�B���u�#$�:���#U�+�	���oo�S���X���]�R��]ѝh8ߣ��OSy{)ey�m�y�����'k�:ˁ���e��8�Sts!�F� ��O���	�BV�c
`w��ǹ�gGrϩ}��1t�&��6l�~8��4A�%��}�.�t��L-2��c~,G_A�if(��	4~NS�M*I���,s�r�����$��.xe���T~+��t:��T��N��T�I��8�'��Px��:WRxeM_�0`�H��b����.���i�7�5�e��L���{�}�M/���� O;�0��M��z�<��K 7m$?ý����^P�7��Da4�h�)݂u�����P:6��e1����lVƦR���)ܭ�Y�7T���S���&e�a�o{�O�@�1R�^�]����_���Ye'�GϿ�%s��0@�[�������<��˅Ǜ=c$~^���G���NE8��w`f7�3!ǄG	X��xًWi�`�w���G��FC��S��S���Kt� �;C�S� cV�{���qb��i����;҃ġF��ǆy�z���
������b�"��Հ0F���j�8,����E��@]�����-S��ktg^5�Qx�L-{qX��N{e�G�$�=P�� �n�(F�[�QQo��2;����J�o<�G?�T��ET�����Y�C������OP�F~�>�8��DsAu����Q��#XÐa����Hw��p�/�ep�/�ũ>��y�;�ojs��`!v�z���]
7z˰��`�ش��q�w�U�b��eh�4�"2���7��ig�3+���\͍�O\����(��[��r�rK�L�:J�D�7DT��/��Л�}�y���˛\���ߍ#�+�ӱ�p��|7[�����X%�9b���Xi��dK1�I&�ҹ0Q�4���6�z5��W��J���u�Ke)��.�ǰh��Q�� V���x�Z�%.�ҋ���N����s�_CW�6`xU2��zB@nq��D��o!  Ŗk�n����~ą��<jWfq�4�^��1��y��>����I��&�ŗ
n�#�OD �\�QF��<�̷�H����Nᜫ��O@����K��2��)��r���1���Uʨ;{@���E�1:�IllF<�t�]�G�6�d8K7DN�`�®[�b�}7�Χ�9��e�N^�?`���o`���Kh����`�1 F�2�������k���2s=��LQ�=� \u�,�:�R6?%C��������Ƿ��1,4�;ں� Q� al�7$׎F̡�q���X@�$2�D[�U���&h�	fh/��v��yB�����f�'�*�a��@���}�Ex=9g�1�7�ݶ15Z4>��Koӹ5�� QU�Aߒp)5�:���b�Ц����I�߱w�4q�j+hqRL���x�Zz�TZ5�X�m�.�����@�u5:�y�"��{��<���u��bXN��ζJ����GF�����1�#�}��~|��I��j�j<��wbw�^D���zD}C�)Ǣ��1Y����zG"0L8b?95��U�gd%,ABxߞ�T�ˮj)�\k3����0���R�O���բ�,78g�m��q5��uO�	���e��i�����I>}`﷙8x�;�L���334��5�-E��,�y3n=WZ5��`ɄWB.�[�����Ό�I\&4�.�u�Tm��1��s�R7Q�Q�䇱{H�M˸qh���P�`����0F�W���h�%��u=���2�����[J�� 8�S^"v��2ܘ��c]��gY�r��3܏q��p�m��C�u���c�����va\��B��6�M&ԅ5�Z�g�˷�鐥����y�rhxW� ުI���$){�Qk�MDW���ڍS#��w��Kw�����}f���ⶂ�)�������zbJ\l}1�ew��Y��c���2�SL�T�2��aT��;�����~0���@�է9hXK���T6����(��D���C^³H�6��Ǝ��Q��)�HЍ݈���n1����B/�������+-�
qoryrm�Y^<1�[	�C˽�D���f�;�Z#�M1�y6B���� �it����`|[���d�^�%p8�vV�h������%��x��^q�����n��b��=����<��i�����v���0R\Rp�AQ�#f4+��֥RQ
,D"1�92�!��2S���ܹ�΃���)�v ޿f���I�=�'�$��B�A����(8P���+�ʁ�<��MO�	7��M��<(�?��%��O%�B'�i��=>�M��GщL�
zc�p���j�`N̚����5�9v��J�>jG$�t�+�*��[B+�@�xZz�^�0Lc����o\ O��]3���~�r#J�'�+D�w��T��QRx�v�S�Ιh.!N=*la#�槂x=��hY"~��g�֊�\�$A_ch�	��))�lmfݕ�Z(:L��NJ|*�Ϟ^^|:
S�DV���p��?49���(���W����(�T6���l�Հt#p�a{�ЁA#�n�BPGQ�CzѸt��A��A5�ot�ԃ�uc�t�/��� �i+��$���_�?P�ܬ��F��b;�Ͽ�y��bs.��ʢ�>q�L���|��鵑σe8�J����ƳqgD0�Mk���x�#���m�o���a�s���M���Vy7}�,"�O> RĤ�XL%)�V<@G���*SBo�e,cZ��1/%1����g4�c;9�����r�O�6ƅ*��>�!��r�mj��Q?�)�>"Eq��u����{G�J����c,�v����z��i�K�21��H��0�41�y��;�T���^@�Ӏ��K�k�f�y҂!����+�f�r7�"/B�ӽuR0� #т�a8�=`n*�[��f5Ӷ�4�"�?'!sp��+4� �~KY�Ȟ��:è���������{�-��G��m�d�,|�%�nV�KD�5T��ʹ0ޓk��:����	�h�σ#)m���b�\��|0(�M�`J�ֻ+
\=i1�+2��,T��8f�M�1��9gaq��_r��eS�H`-�,YX�.�I�\�[m���/�yB΁1~oϛZ~	�x<�Q��	ͺZ�l�]�j6�7ѹ��",���w�$���� <��(���֐6�!l� ���n9�\Ac����|�."����ֶ�*��_j7�uJ���x��kGT�$k]'�^ץ�ĕǠ�XG�����$$LF`���~Qg���ج7�w.�#�)��O���!7�El����䮕Z<e^�7E%"�!"�'O�^�6�mHq�?��۹I��A�辂���PC����?״���a�7�e�^�ʀ�~�#Lea�����
���M��=��[dƦ.+�XY%q��Iܤ d=(���i�\�نy�(��Ά�����Tv8;P��&G��40h� �GI���C���1'��I�֩�c���t�	����^��{4�$�,.��D�>�zA���<� �<;�Y��E{F��/�����2�lhIs�61l��4��{[.R
�Ŕ?scW�.I�*��w�܈�I҃���jR ��P���őݨ�4�V�?E2��X����`9��I����Zt�N�
I_��T�
O��bhDLT�{� ۹��1 D�����ƌ�4tĖ!�xf5��P�əA��"��j�)^��L���8j��Y��Hd�[����~S��Q���+����DK-3�͈�+Z <mr�񳗠�|��V�j�ڤ�q�� �x>C�����I?���+�n,��:YF4�KZxhh5����'ޟ�?�C��������O���Ȃ�9�{V�cQ���՜F���i2=> b/3�=<�q�ة"�`���H�W���3��.=�O�������])�j�Κqu�N
�����5��T�<��N�gC�X.鞳'�͒��t�
�!y������/�w����IN���랩ɩ��� ���X��ii�ğ��.EY�����d�%t@��')�ڰ��g�v�qdػ���-����8���	]����xY`�ϧ�<�]_b��1>1�<V]�3��cv����_�ƾ��j�V'�W��̵FP�1;�Ju����hI�!�"(ޢ9�VzAS�Wcm�7FA����cN�,�cȴ&��"x���M�*��2�j>���o�0�5G0�=ԩ� �,,���8��L7�
�W����I�0��W=N��&A�>�Y��=�<D�1�0�4L�pף��]�+S+�٧nØ�i��ѣ����ke�R�;��	hȊG�<}�2Ϭg߉yi}?|W�gG�w����R{����j�����%�݆9;GD�����K���R0]�Kh�\��S�H�%��I/(Ǻ5&2�	I����o?���c�q���������>�eOi��yZ�*ܭM�� �$� ��jS�۪����X���;�ET�Bӕ�T8&߶�+�L��	��[�F!�� ��~0�vE�	L8\z|_c R�����z���QZeH��{U$wfU읪.k(��h�߲��Ȑ �&�Q�z3�T�|�G�Hr��;:'D U�x��? � �R"�����6\�ħF5a�N#�9ł�i��:n�%z\����{����`�8�e wu�0���>�S7��=@���g�oC�C�iv��py6!�^[��uq}�JZ�)�����;Q�NsH����5���u�~�A��Klf�	P��w{���6�f��5H�ix�ޭ,���,X��N�u��3X�&>����I儔�{6z0��Ɂ�ܟ�7�qBG��6E��<�� �I��YW�'kD3�^�,y�ߒ���q�{�����l9v1�K��~�pb6�,�n4?���(Þ%���G#7�m�ȶtV��3�{fN�e�+�*~�Î�Q }��E1��'i��DD��U�?�,j|��c��5#�΂��j%�~#�*o�ʞ��Wl�Q1���"����T�q;��KN�B�[E�T�Gć��xx�p ݸ���Ζ{anQ�b�߷���^�Wd��gtY�ue.�g*i�������e��x�X���JX���ʡ��" �nYQr]����5��_ k���3�k�Bqv�nbOϐ�"Z���ڕ�50V���9��|Q���za�m�Z����y9=��L��Z}���|���f���qrWT��!����wc(H?>Le*�dvGK������P�َ/̥v$�*@�'u��"������V��`W�5�m�z쒜Y";is��S��>�.cd�@��>s�F9���+�!�pEiMr&DB9�!�$ڼ�IԻЅ����wk��?����׊�6WI�e�6�{&&�t�J����f�%�,��:Cg:�'�u���T�~%����G*q��<���5�m�_J����:4菮��l��"��R��Rg�*_��ʯl{b�J�����?|��'N��af�:�縓������"a�L��"����y��u�JB��T��<f�����#E�l���ޟJ�@
�����ޞ���gB��Xo�~���*]��o:%�Д�-�S���Bo5x{rN��\��H;S��j��'�AGF�w�O$�� _�U�㶸:e�6�OZ�dcӍ�);�$���Ȓa�q����q��uo� ����#A�ӲQU��-�y9$(�3t�lw��r�|Y{�;H#�4��zn���dB����m|���d՜��#��e).���+ٰ����J�߾c�4��UACД
�p(����MҜ��O�ｹy
�C�hři»UI<#����.�zb���s�S�Z��^�7�29�m�Y�x�W���9�U�V4Bt�L8�ff�袶����e?K
��b�{n��A)W0>-V^�d��n�?�$��H��~�.�`'���bDx'��J5/^��2m�L��� ]�/܈_��&�����2��p�n7I:��6X7��GA�;��0�;��`�%$%���kX�����(�m����5���Y:��d��#x�]���y��#1���QOD�]�d]'Nt��y�K9�y�^��_�mq�d ��C�J����K,7��t���T��[h¨*OzW3�9=�~��L
��N���ߊ�R�����>��	�f��qwt���v�B�~V1j^��XȦ��9K�Lm���B�G&��,�ֈ��!g�"^�<&%:�츠ȃ�)�F�c!�{h�#�o)�g�!͆�|``���e��t
G׹��@��="���LG���S�;��孭AmV3��E
�U������z<���*���b����z"H�K��g�Ǒ���7H�ѱ?V��CjvH-p�|��>ޚV`u�ņ�&#_3��o�5��c2��W\f��	'���]��'��y� }cA��U�mC�<EA��| ��DJ�YT��q�� }��	�E�2����� ZC�Nz>V �!.Y3�q".9:��&���g��&��+z���S6�&t��"��Q�f�o ���r�-y�n�+��,i�.W�_/���S��8.��Փ��%�[Rk��d4��-�A�u^-'�Wv��&8���#J�����mpաz�C��SH!�(S/p�`����~#����
�	����[xp��4�~%�B�m�c</�(D�ɭE��5��Kh}�ֆQ�?�yn+�\��	�� �k����i��2q�
���`F"�#НR���]kx�	&̀uR��wv���a��Ց6��T�@�Ÿp����'����D9d|�#��&ݙ�sT�N.l4WEQY�Z.g�wD!��@���6[�u�� �޵�f�Qτ�9�A�TuG�}��:H�_	�K��]�$˼!�<�#N�dR$K����!j ,6�ѯ��V�]�V���B�KK[��c�x̩Io���V,��Չ8�"�UE|�BZ��t �D� P"
��T%$�7<ɔ�`��x���ꬺV�vs�l4y��BM	��K����~��0�����g�����>_W�5�7&8�����Х�W�XU�+Yr#�䲖������x�4��l���|e?� ,m.������4�<2��ueY�l�..��t ���׆Y\K<��-�FhmB�o8]������Q�fO����n9��6�]��@YEN_l&��2��&N�����ڨ%���BJC?�G�����Zd��(�C��Ǒ/�{�[��823~���������|w���X�؀�3�}}���|���Y�h0k�`�&����C�$�A��=�Gp� ��\��U�F��L�K7�P����A�p���QVlha�Sg*lW��(ǴB@����UT���8+;J,�.�k:`/�G��8�x�k��>ZH(�!�ד�������UZ�O�-��:/ݺ!~�Lʽۚ��L�oՋ�K� xJO+?�N\����������;t�[ޜa(������~���k���/�#0�l.ώ^��W��DU<����-Td�ş7���1t�d���yݴ�L��]����|��7��N�Y���W9)د���,$�b�CFT`� � �l����^dv�)w�P�j�W>,sW�g�	~����C*�_=
g�P��#��.zY�}��t�)ç<>��� ������_M%J��\�~J��{
suk:���{1\��������0�tq��-Pl%�y�P�ȏ�^@���n��Z�����,i�3gRװev�0�X�g�H����"�¶��V.�y[)����2i;B*H:WH�ÊD�ܫ��WԓƳ�[|9@`^Ӽ��t@��u��?��9\~�������,:�Y�k~t ���R�Δ�o��A����n!��^��~,���?w�Z z�f�r�[�Yl~(l�D�S�������1��-S�Ƕ��=޼=Y=�^�$t�א�P%S9<�dn����o�r��#�-�)�\vg(d���rQ��U���]C�+l~C���)Q����xf��.m �C�l|8�3 ?��ݤ1�-���J��Q\ڦ'ϡ���pZX�26
���ʟ�u=O`�Yr>�������f��fT��#�T�(����~��:௷���/hf�e�*LH��;���d��� Z�o�-�+�NG���+��c���Jf�#����F)�q)}���c�_fr��"-�6b�2p�p���)�#��~���9�����Fp�����E��]w�(�o������Mǯ���I�lEø,u�w���%�-�飦mEِ���!�+[6O%Y��7�[��)o���E����;.)P�}"Ug��]�	
����^M���X�|qN�ݘ���U�]��Ʌ��������^�H��~5�#ɏ>����x1�TN��X���V�7W�S�&b﷿��%���	^���7��*�(�B�Rl�T�Ԝ�z�tO��!H4��q�ʹ�6IИ;RPl�s�0 ɼ�����)�(]b$���8]�#�@j�e�TC�7�x5<{r��Y�5���@�n��
�yFv#��W-'�������P�Ѝ�jb�RSk��.���,,S�$T	����p8	;e��c��j>Hef��>!���n�Yb�8,v#�@�.�~۷Ku��>��d�n������>\������[��j��k�`
����аY�6]8��c>^U�5�BI�����uQ~������?fZj���j�<"!kB3�b|�� �(�� [%a*�1�"S�wnQ���Q5&L��w�|$���DwV�A�n��Rv�y25`g��~�3�2%��1������Ǐ��d���t�~g���?�ev[>3P؃��[]?}Ч����r� :.�9��ԥ���8��z��ċ/�gF�<�	�5&�|k�D#�>�Ⱦ���E�Y�Ud�'@A�G�E�����]'�3���`ea�%K��V�������Q����~Df�Ϥ��z0Z9�c�
��4�O��L0Q�G������R;��j��$��q��<) �����iG�վ��M^�/�9y�x4R���c���x�Q҄]_\�d�ϨpX���a��+�֣��E�A(��6��k��=�y޳�t���m����N��ּ��Zt4$p�x��Y�ԧ?�i��\B�wV���D��A�MX�~�uG{�k�P�F������ ����ĻM�A'J(���Ć�1�7�Yԍ��D[�fði�s�&1jB��`^Z�(-*i\J��[�m�-��q�p`fb�e�g��)ň���NP$��Mq�r�y"�jT➤�~s��<~�>\ �F��%�=�HdѨ�I	�V_%l2%!�4.a�����[������|��?���]��U��|��X�*
�Ih�%wy�2B���������N6~����I����l�Oc���kQ]��؟h$'��D&����u[������}Hc�Ud���	 �0����*��b�=�)a��cm���[Q�yY��ZHL���|�AA;��Ē�t����'�ф[w��� �wY^��C��
�&�RIm�ʉ�##ѫ�=T>Z"�o�ŗ���-p������%$$dNNb��`|��i��]���i�}�7�4�����!�t�$�1Y*�hK����~�g�����<����a������x5_:7{�˱ȝXa���M���ރ	�¨��Qi�s�Ӓ��,%ϒ�au�FKj�P:� 8��IQ�ٮ�I��H~H�����%�;�s�"�*5����e�껌����Rռ,�.��Dt�4��^Z��>i1&Z�U�h�>Ԭ�&�8�ɴ���5�D���sc(8d�PZՙ����ؾ�˂�V ¹j.�'1��z]H۟�N	���T�2J��3;�����m&�Us(ӊ͛��5 �~����� �kY� ��s��I1Җ'���(0����i�a��G{�[u���-A�3ZݙJ{+���Y�����Ђ�r�WF"	�rR�޻��*�b_�"��F���9h+s�-7�>�Z�G�d���������Ƴ�O�Ӷ3H*D��`n�[�{��3����f��b%��<�x�Aְ�v�=j��"���ǡl�,�;��_�:-�l;H�T�_IC~�O�ݒ�W��)/�ċ��R�F���K��A�PIGm}ԅE��L�p-���(ᓞ�l`����Rk���� gݲHڷ������C�����Ȟ.�p���`d�Y��kkpn��M�d�6�J�L>ʚ� �!,V�4p�9�Ρ�<�&�cɒ-�D*u}���r��"����ͩ�,�y��?:EG��-ݫ�N7���1جq#Q��>%�*}|(Lɷ��++�-�����&�� �� h#j
'��P�n�y(W0	�TDQL=�ō���)bS�h�RE?O���b��%{=�4ndI�� ����:�����n�`UO�̻v-���#�y_S�(1�ʈO'5�*�ha�Z��
��u�ݍx�8�y�{�Z�g��s3�\e�I�y�c�nr�V!�C��<��M�M��̵�@f�mp�C��x�����Tn`/B���.���#���`ܹK_�� [is2*76�%�1��?��g(�p���&T{}�D��6Sⴾ���
���=N��`Ow]�LL�����|o�HP�<�`Q0��]�.?��E���h��%$Y-��t0Y^z@)rK���٪��9�A��B����g]q�sW"��v�C�-�i+�V��"���<�TM�!��;L���m�=7a�+XE�J:�}"��>P�o_�܌zFxӃwjq~7��YZ*j�Ă������T��܌]����jd6o� �r�x2���H�o(�
����.�d����=5�(bp�3�y2��n��R
�
�%��l������(��īuR�-4�+2��㥇2�g���v�&���͓��$��"��%�uP���d��:*r{�u� ���J�qc�=�Ad��-�e�j�e|:��O,z��חz�NI��ż�G���}3�h�J���J�"��	�*,Ϭv�	��̌���ԇ�v$�K��&�㪩4YR��jliQ��c`�N�� ��c���
D�~**���(���*o�TI�]��Sc
��W$[N���҂�5o�����|<���il�f��q�l ���V��[�����O�?�%��	�*"�L���H�Ɏ���~|�J+U?j��3���ca�1�na�Ͽ�&L����h�F�z�����!�Ӻ����R��:ފ�����:�,`j"casp��,��ed�$�~i��j8:ۯ�q�o�!��ENlf�t�@ŁZ�i���OD7�.��.�������p.F�3/*#'R95!��� ܂��\$�W��p��N��g]G��|�/���\I�� e�
C��u�1�dB�<ze�~�/��}93�U,��I�_s��s@n�t�V���^��D�V� �B���t�*᪍�q�{�L[�C��;J����q�%��l�)�EP�5���]�ȱG+�x�������,Q�p�b�Ǌq*�+��G.�u��������V��x�'Ái/+ʒ��x[�q\�l�ke�f5�Li>������Hv=(�o`�^'�0�}�*6n�9��+�$����i�'3�Q"�P��B7~�CIN-D6�)�]>�@�L�QI�?$��Ӳ���eB��L�({�7v'5n����<��l~лu\;8W����#�r���_�d�t�ɉ6�r�qVR�J>�V�t��#���SJ;ɍ�K�kZ_"�G:�o/������q�b9�&�.�AkN��dB^	���5}��0[�U�;ܣP�M�Wo�\���V���6�^C��Q
�m��9 H�I=P���T^���|���j⻅�t��
v��w<Fd�?Z���~-X�&F`�řmS����58�"�#Ҥ�ַ9��֎A���H�{�0�Ƅ��m(PM7h\F[�DB#�����#w��q_��Q��H��E���T��}�����l��-���2��s���� p�P��Ҿa���c90+���U�uy�1��m�hjEW���ɸ�/��p��v�S����=O�8�� t��K_@C�J�he���-�88�G���.�&;Igzm5z�����jtz����{� ���}��rHsE[
���>����^j��s�4)�������:HR���.5�3GTwt�]U�k����SK��rzW8 8u�\��:;�oQ��sz�)bӎ%Ƥ���ͭ`�K�Z�IV�)@;���H\tg�~Rp�0�YY��[�,�Ē3hgo�E_zvY. 6d�Y;d���y�Zkvx�A��x;mS!A�&\�E�`	���:o�r� |�?s~�����6��l��[��Wy�*h��y,��[RÁ
�7!�{� �𽁵��mS5�P���*2���DB����,�.؏���~�1�Gj�P���[�� �NW�����}�;W���ob�ޔKh#����1�j�4SIzX����` ��픫�e<03}�I5��0�er�e" ���/0��6t�K˚���m�!�v�i*�un���v��!��iB�4�R��ڌx��I{�g��?�Yi]�1�y�����bwٻ md�<i���A���ؔ���b3�y\n��8rh�t�B	3�H�P��5/L1%݈=Ȝ?��}W1��dj�n�'6�y���w��^�$ic?K�Ȋ��;o��vNxd�����V���բ8Alj/�V���"���X�R`|������v}B�{ǔՃ�t=vO�$qԲ��a���
�<`�"�������05���޾�f��� ?��>wʋ#���粳Z����c�y�y2Ck��hQ۹�}���}}b�aQ��Ŷ[X1Ġ�ڰ�	�Ȃp6}�eMa,�[S���?P�W��_��`���0��A�jfĲ�;)|�r��m�"���/t��¢p���9[AiB��_<s�9(��5��Yc��������]*�Y��f��4h�u/�"BA�Wl��#��s��g�Tl6"�Xv.T�U���W����޿?hFP �D~'8נ��/\ק�]gN%�}�\����H=0�[ �[��2#Z��� �tuc�Ê���u�:읉߻a����������(���itl�Ѽ-4�ZS��=N2���b�8?��h��A��C
��j7�A�=�4Dܢ�eq P׈�RiBD_���v��FyE±Ņƞ��L̈�)�����������_��-՝:�1 ��L�FTZ$l�B��I�
�.���i��_�3�Uy�qgU�N���m�>M�������ov��4��n����sF�AHU���k(��eX��<��qJQ��a��g�6�����w[Þ+U�/ֲ��.ڂ��Z�l��kD �Ƀ���:���x1A�L6]�;�ƦD��)⹄8~��Oa�2���z:�t:�bw�Q��Ϊ���������$�2�fHS0�l��i����w>&��o6����0�FZ!�7b�o��3��%Tn��	#�޲[�S]S;a�ϲ'V����=�5��l6�`"�㾇�UiK3�����Y�ZP�aw�\�����(�E� ����j#X4S2��&�D�=���uL���?;����=%�8�R��ǷE�P�@�G�w���~w�SQ�yjA�A�`���c6ΛL?��7y�"
�	f�1��^����^2��P���ի�͆Y��MuI�}C�pr��A��
����h����S��"?���~��n�bIr��;�a��R��Ͱ��]픗,-�e �#�M]vky�ı�&7\�x���=�,	����"�<
�e����cl �9ޭ��5���U� �8�y^v�re��:v�����A���,��ǄCҦ���B��@2ʂ��jO���6/�U�N��� |����O� ��P'�q�\���Dy&�T��s�6���TK�u�.��dJ�_��␫G���*�}5|���c�m5���xV9�˟ h�A�v�#A�z�P�4R!���8r�;�=��s�jy�2	G�L��r�{�=�0�*J�Bj.�Y��Ju�be����P�I�\_��.X���L���u��e�ӓ���]c�
�z̳���XC��d݉&������Hq�;����u�]�sƞz���� ~�AjEHb�4��1�n��Sq��ƽ'��fp���XRӪ'��#��	�c��q)tx�Ok�z¤ק�)�X`�Q�� ��F�vu>��]'����id!3D�Ը�	6	&����.p*�,�㎬�MΛ�al������P?=9�<ɷ��>J�8�S�z��xP�Rch�H󌩊?:I5�^�'Ddr�8�<JՓ�E�q���� /�U\�L0���W/*2	���.�t�A<t�2d���_��-(rW�y��؋:*H��������v`+D]�X�Mi�f�f,)��3w�;n`q�0��m͝fq����Vm2uJ�h4�r�W���c�aQ�,Й��%����b R4����SwP���NΘ�A���F%�g��p�����E��Ăܸq��yP;��K�����R�zXv�qo?�)�4���݉m�c�	h�/�&d�y�zz4�$�#D7_�.�0L�8�� �~8ZO���4c��֞�!YR�d���l�<1�$�al_ٺ��&�
��s�@�Fŧc���@l������ﳻ�]��Ğ�Y|�ڏ�tg��_P�k�Ç֞��]�e�G�w`?9Z|��Gxƚ.��M[��gf��Yj�z���Dt/�����ΣS��ۨ$�K�����8�A���WWnj��	HĴt:e�����* �u��l���?W��8�=��}:"ۼ�a�C54���W��ӈ��`v�p��ۯ�~2�#�K۸���̋?$���9���m��-�5�!�\��DY�����S���̚�G�Qt��T�wU:��r�p�F�]��� ���M�vޑ/�`�m>��C��GyK]9LX�_M9C� aњ�I�6B֍��.�e)�[�u�wڝ�L�J{��Ǥ����6��*���.d�d��4{`�>��}W;�+��1s
am+ڌ,^����sMQCR�{j���tK��9��M�] ų�@��L��{Ie�P�Ybg���<�!�ֳm>m#��8��)6���b>J�鳒6�K0�Zq�m��3��Q�C����."����S����g���M�X�P?~R6s���p�򠽭�9��������iaMbMQ�Fg�'� �q�Ν�^%~�|Z%��{?���l�Q��ب�X(�J}����`e��Q�CƠ��w�y-_�0�՚��
����0�Zj7���^����4q�_�&�����N� %5-�8I����N+S��.��/�ʜ�������HV��c|H��IP�j �$�������*f��Dh%.�2&-�$Y����#{[͸	VyO�-��<bm��U�(�7����d����7����|h����g�공p��գp��Z(=J���C���l����2�� +�P^q������wo���1�kf�N�2|3j���g��.3��~nEgq?+p��r��>����C���Gbɋ�	���TkM�~鑋�����x����q��/_��="������M�Z����(�W�����V(^E�;��V�b��Lq�eg=�J+e*,�����q�N4�À���~d�,��fU�����j��FT:�i�TP�ԙ2�(�����~���)r,������l�/����[���^����̓�X�qP��f�Rj�ku�I(zY�9k�K��S��6NO���Q�ky\�
A6tu�
�>0�$�`��@��#��v����57ż��9Y`2߳�𐙓�)l݄-2@�M�&O���=�״��6ĺ�q��SM��I��Oi9����!���P���=
~��~ �:�iG�rK ���X���tE	�o���B[�{Vu��C�6��k%d�s�_&/QO�$��nC��z H]h/R���1��͟,��=:�y�!�E�֯�fV	l-u ��}������w�g"׿��h�̕X� u\2��%`�O�ki�'B'��F��G���b͑�y�bA�_7��˽Х�ƑW�u	�ˊn�-�	�ҟn�Άؔ)(�~/��j�م 
�,I�h3�g��E�Q��;0�)��[Dj������
4�	Lv���сl1@�/G'$
ӆ�n�Dy���TY�Dh�A6ᅜ�G�V�i��&L�����kO)��?]�kX^nɉ�FW{8�9(���X�[Z+���AS��t �ئ��dpiK�]�&�VIӍ@�^���g���îH�*�N�!)#C�����L_��q��\��X�����^�Ά�PӬfS��7���.Z�0�8�"k�,k��-�>r���K���:����C_U�)w�u��C�AZs'�8����@�%=
C2��'w��/$(��5�tD�"q������;�)N- N���bR�~Z�z���8W���\���0����)k�14�-T����h��F�����GD^��x1 �M!���AT�B���E��#(q�*��i�^�2���A=�G���}iO�`}x��R��~4̉�^N��&C��_�������Y�̾��O4Ƀ����i�n8�]B�n}��p���Ҋg[F5y}�z�ؒ/]���"����V�B�N߬R��"ί��#�%u�>��%d�״=���}�V�2U�U�8m�S���*��Ŋ|~6q�wWOD�����uT������8$�"� \:��`}%�n��� ��&g�N�E�><Q���B�J��%�v6ЈIa�-�p���s��l�TFJy��<�-p�u8�M�BڵD~�������q��IjY\�������x�Ԙ G�1�J4�]}���4���?:�F��ԍұ�c�9��88Hl�3�gL���n6���Hλ�$8U�� ��"]�#"�?q���́�NAȭZ����GT�����}�p>���+�p�7���4(w���	�̹��*���S?�s��r�:��KaL�<8�d&�B0�6-�m�����*Q�l��5�o�^�o:�e�H=f�ih#,2�x�p	�Isv�/��802E�]�u�/������1��@?-K/���A��*�7iz/o�}h���[|��r�G}@�,�p
���7��v�;嘟j͞bP��!Sd!�����BK�׹��/qx�0�r?R�eo|�U��[��	�ďb�a�<���NZ׭�C�ќmE��l$@��7����e'J�>�@��b�K2�Rc�H��@��f]Ȇ��Y�6����`+�=(u�����u�Q��8�7(������ P�]�ARD�=�Y�/�a��(D��C ��Q�-X	���B(_6}G~Ex$�E��-��;�"�(�4(	��vWH`�<�C\`X�q���kA�~�Z���P^G��x�J��_F�� ��g������b>�.��8�{�䬰������m
Ӧ5����R1��=B����%���F�{�2�`ȃ{t���!N8����X��H�w�؟[�|��͆s[+bd�'��2
fE@Ǧ��g��o�P���lx8�6~�{�#6R\D T�iv~�;b��V�]<d�� ��<�r���1	ΉX��5�Q�$�� �	)T��Ö�.+�{F���W��v�j	9*(���c[*�׺�b�O��SRĭ�*�������h��a����80�_m{��t������▊���b!� ��������y���W9~�?�]��!�Tr�)��?A<XvYל����QU%�X=����6�C��A)J�O�w8߉L��Q�Fd��naS5v���w�Z����/Ӿ��ӿI�����