��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����xLM�����`,5?p�"���N��}߳�^'��v�Y|'�XR��f����mM�x�p�xV#ڇ��76{��)����L���h�:��+A���9ߨ-� rā�SZ )����C.��&0C]�-��[�3�-���+��պݣ�k�J�vo`�A�����f����u�X���v�=�а���]Q�Wۿ�߸�=_Q�X����j>��Zw�K��SvX��ƥ.���#�����Z�0���#7{��\S$��@1I�QX~TQ�E��db����۰� ���>0�%�9�j汈��}��1� ��2���h�G��SeY�a���	'<x�p��k�H`�H�j^y�0�s�78+���ֳ�`�R3dW��_��{p[�?$�s0��#�zS�_��bH
�c�p�IL7]� |����Q�� ��Rr���=��E즕2%�����`�^��l�q-�]�p��jf��Ӽ-f%H���ȳ�>��+���M�71��4_�) 3�46h�rb�J�W� k�h~K0�>P$�_n)���5�r�j��W�J&޴o��$>��6��ŀ�;A~<6P��K�~��f��*I
�Z��}`q���ApC��n���g���3��-�іrO�mF���,�$��@�BI�q�}��Ȥ֐����î�䂧��@������U���vU������ �T#K@f�㯁����|95<@���+�-�)�����K���FI�k���*@�m&���
���ma1[�2�u�I�\�U�yu���o�|��2����;�W�W�}P�K>%5�'�8���׫=����k��,�t�M�0�8]q3���N���GvZ�i�+ C�e
��Ќ�S�v<%���q��e_��
�k�夞��>ZO7E~��5k�TW Aod��eE���G���ɑ-'���?�G$����ќ����8ɸ+ 5ʗ���l�d��,�J�
�^�3b,�����J����#n�zK����z�&��;|�\�^���'e�W�����">�w*	FO�Δ��v�ƺ����U�
��Gg�Ʃ����b�7U�/M�T�}����g��40@���f�������Bڿ6t�1["��rI<�(�d�LE@"��#"`����Aզ�Ů���(F�q�}��LI�q>#�fHֈ�K����/�h�<���7P��x�����,Bis�s�F�
K�bTlR��z�4X�kG��`m�sII�5�E
^H�!]싴�F�v�{��O��j&ef��r=�D֢W��_���s��f�|f2��B�cAI�@:�ݾ�9+C{^m��g"���)p����&V����a\�����v�	�'��
�Jd��-��}�5����.#�|�B]�!��Ǡ��������ZsǮ�-ڧa7���7������9���M�r�mN-e����:°���I�T�X#]�-ѳL�M������o.I�n(��P-O��P,�>7n����$�>��B>�c"��|s#�S6�y~
��p�A�)�7ΐ���� �k�۩�1N9�Xh͡��ñ�#1��^�U���k�;mz�i4�UB��yř���w�YTut%ᗆNj�����Tn�C'1c��e���vE��>_�~Oq�a	��m��Ol�N��ppT
�L�C,�n"fG�D��F��B�$����J�f�g�Cy8�q�i����:N��v�S.K����P� �}��;���&�h,p�Ti^w�b	��'�0��R�ԫ$?�C=Od�7MujLړ���F�PV����WPh��u30A��m;�1����_Pٹ
��s�扚��9��X�F�\+A�bW��1��	t��-�,�o��ě�s{�O����Gߙ?�{�̳e�gµ��EQ1>��O��� �@�&��������z�ƥ8�#I���)�i��l����8>��r�v\���v�� j��X~D��H���|ݣ¦"���p-͖���������:z�����xH�"I��ZdD)�CTs^�Q$�
R��hzv��%�ޔ>���g͔JY`�=wUӨsoʃ��;)�yW)Q����B[*�r	7WW�R����B  ��T.����	��S>�$i}��S���Xh�@oF�?�r��ƴ�q/!�M�����"��qѹ�]/묲�A���y�k�U�L���0gvƨ�S!�?ü�'^��xp�{�����Ӝܔ
S6 lu.`ꇪD� hr��ek}�S�xTn[R�7��0ĺɶd��n�6��5в�f��خ��<�ݜiD把 �}�o��&��Op�}V�i�!�Pn�2����s���O�GR�l!���e!<�Vƅ/�+hl��C�8� ���&��:�%���?��F�K&|_�e�3h4廏��>뒭��ۤOi�Mx^��
�i39�V��h�S.��^��Нk�#�F�,U�0G�%͎��os�Q3�^����m�jC����"���m0�\㮘�Bh[TRoݑߞ����%�S'G��Уׅ�j���u�v�VT�\ hǳ)�D$�����)��/�[:z���~mb�@��S�W4�y�:nb�x�2�re����̑�W�Q��K�������y�Sq�k IM���ȉ��ၿG9�*���h�7A䅻cW;�����V�D�Xh�՝J�X�*ue0=���k��v2ǋ��0�G���m�n�������mE#ݣ�g�g���|I�:�l9g�K8H5�C��� ������ Vq�9c��b�O�w�-�8���RJ���,�����2��w�ik'_s���2/C���(+L}v91LBur�卲l
�}V�7���L��:0�Q�l��qk�!#V����c�Oqg,�p�Ww͛�~�/��{%O�L�+~5���.��+�k�^�\̭0Bk��ֺx^��eԚT�Ű��	�~CX�p�E��W��uu|+�n�͠GEVf'��)ز �}EҤC�`�&��1  ��'<|=���h���y���'�hE�h8��MB$�ձg�H�e,�`㉰qJ@'��+��R�Ț%Aw �|3����駹d��i���{7N
�E�8��~Lb��J�  %� /^dw��Kο��h�ڹ����qn�$����� PB䫲+�&�8YT�Ӯ�LU��&�nKk�Ho�P��!8a�-��,9P��!!��mK���<� �נU������]�y�
!�S�,pL��������C8�渖�W�gM�/Tcx�Y���nk�}��D��=���������[�V��p���{�d�w�<�6Ӑh�'���cV��f �F��I$T�5��?ZnzL��A��r꧝aE�I/�|t���ڠ	�&I�2���vd×h!��	��[���7e��a��b��n��0������iL���-ћ����c�{�h��\��I��H�;0��l_�#�#p[�Y�u�\Kd�G�kAv�H��9�0�/��r�]k;���U=���`��j[�/��	������?#9-Պ\��i��rj���	7Fe��=#"�eW@��ŧ�D5���Dٽ�m����<3��:��#Ϳ�âmf��7<~r�6}�$�:��x�Xt]����6b�?��dg
�Hq-�s���*�/<�b:V�%ٽ���D�ܐE��"�Y�b ���H
$�L�֊���Y���v4ڼ�.�:Uqu$4A�;vx$�B�Xw�5���<�j�d� *	*E����{�߶L���}�ᢜ��D��VA��/�sq5����A�N�{n���l�/[]��q�Kq ��gO@�k�dIBО����,�_����zfR�`�Wܔ���W��GF����ws�L��%UUc� ��)_&��w�Ґ��E���ejAWg�8H�͙��, �+bX�_H����g�S�Sh�`�{��{ף��I\	���6��H�I�"�U$dd�@;�����SA^!V�1n��(V�r{(JP=��5^�:X�xO[F��}�Rx0��O��S9��Xl�v=�B�S��# �nuS�VU��0<(�2����mp�s{9Qy�Z&�KLT�Ȥ�dV��/%�wA�b@�uk�ʚ
D0�pb�0�p&[@��H��n\����m�:�i��Ɉ�?j�H	5�ü%�X��
7���I�"�I�Շe4��y2S������IijlC�G+J!�6u�g�N�U��Z��^U�T����\f��Z��z��	4�������P�2��B��]����k� �A�c�<h�U��SJmD���$��t�R�<2�d%2s��*���Hz6S�:�=��d-!�����
���\��i���St���D��D�Z����4)�>��y�'l��jm�~ܧ�]�&r�["����d8���~�OȎ϶���-���
@FtP�as����RJ���\+�����i�0�e����&D���l�!)����;AWM2�.)����צF�d�7�7=�S������Ky���nQ�%G��}V�`�<KU�g�W[8��3c��������L<����-���Q��<�p�X�u��RR�F$�;��1��"Rf��y�A:U�����!H��_�,��@���̷�7� �5��2Z�Ҷ�C��B � �0U��v{w®�
"R���(�����V��w�<�Pc?k�"(���+O:�:��|��w{4[Z�^{G~�[J��r��J�qq�5�O�L����+R�y2�y��j`� :A��8C��P��6qz�ҀG�I>�M��4<A�	@ZV�G�2?}���0�z	�yY�}�`h�?�8&�K��f�\�-9��J��]�9�w�#�c�(f+�QWy"�"}��&/�W.2� o�T��*VصX��jl��	���	���
H�HVz��D
!�E��$q���2-�N����i��hM��@+r�j�D�I6a�&`c�ɠhR̡�%W�/a� ��)k�!��lYE�	/�[��l�
��+�5Q��� �����sng��������P����'�S�"f��ӊ�Q���\��LI���V�������� [M��U�w-��,7K�/S�Q"cf=�x��.q�{m*�F<�C��ћ�c���_�whN��C�P�Z��Z�-��ן�%s*5>�2��̋�J=3���(��#��Ǝ0�E�?�iId� ��u�ģ�6�E����W�U�ף~C(*`��I?���JI�٨�˷3�w3-|f�݉��	Q�6��Q/,4x�*���5,�9�źf�t�qx
�$r�Nn:(s&�&��>��n� k y�����!2���2�C2�5rM���(z����$��v���`RĀ�S�{8�@W�wy8߲H�v�*�����V�7��O�1?˂Y���6Hv���x�ǲ��Oy'�r�D�/�i�3�_��F\8`��}D�-;��ofQ��l�2ݼN���y2$��+`������{%!x�t���`����ADN���q�j��f�Z��ysg��ul�/�����B�ll8U}�[��c���I��`��Pk�O_z��iW���ؗe��y�΍�#E��P�0��.�� -S�'�i~|0�{u7v��KU0�;����YX���8�0�>MV�Q��Io`L[?����}.�Vj��]X� i�L�ꂃ�y������]I���~���4"�bk笤�春3���Zk>�	2���u�L��I�k�u7)ޟXt(Ԃ��_~��b/�QX��s�Q)��!A�R"+�kβo�&gB[l��U�V@�-`�u��0v��Ū=�y��؏�4�)"�g�m�0 Q�(����
�J��>�F�l�t�!m:N�
c:�:��s_���{r�K�'���[efT�>�2�qo).e� ���񲵖��;�lF�c0���`|�%U��,��&��9���l���w�W{��sd<B$��X�V$���"��v�L����
?����l��@s)c*�x#83�Ƽ��ؠ$����2�7����� ܛX���qq�� ��Y���o���$68s�3-ǧ�@�Qj�]2�$u�#j2��h}��y*?H͒Z�ZGݤ��#�
�7�L�Ҡ��:5��l��8�!��3���o����i/p����]���?�p�GÓI��ё�sl�	�y�S��cX=���ԺL��6���1�9���|��o�#4(�Bv"��XZ�`&ś۫����@�Y$����~�>�dЉ��C��W��o̉}��Em���b��x'~g����;�vd��YQW4c��:HĲSީ��<`�/�9�[��2��ձ*��-��w�xʴ�m�r��ׅ�2�'�o�e
��
�;�RS�mض�q��	��D��ׂP�.�MJ�ս���B1�x�����5�Ge�I�k���[X�����.��r���"��+��:p�����ó���f���Q00)Y�!g�
�a��h�f���_Ռ�n�W��z���S�)ս�=��O��@�V^��`�>b��#�v���ۇ%���|^n�;2OX{4әf�Ie:�Mل�)�c$���689ia���M��5��ݲyv�N���h/�
���~<���*�W�i��4x��m1����'���Ö����1�g"�ͯ%�R8/��	��m;�:�R�?���8���V�ԫR�-�)���u�*y�@}�I�(c���X|5l���|��%��eO̊�_toΞ�F"��m߃k���>S�φJ���%pV��w8�Ќ�
���T���2%���ï� F�2�I�}�
��B��>=WG��o�@7*ޮUN��}/u�,�6��E�6��0 w�������Q<�\6z��a`z�#��q}�4j_IH/�$�$�R���״nn0C_.q*$F[�: ^�ϣ� D)K�K����Qb�aNaoö�,���^��k�Ϻ�@�u2��V6�nu�������^v�4�H��LF\?&5D�Q�ڶ�L���Z1NV�i�����6}��C��%9R,�����AW�W��$��r���iBg�P!�tU�_���V��Gʓ^o���Q0�[�|����'K
��lt���!�ifj��a�
�ۚU�n����	r�3�:ֻ$� e�t�1��R
*������8�@�K�P*z'* ߍ.���*xu<w�]��YN/U���i?6׿`mՆ_%�:JM�����W�08o�q��hs���]�����ܸ�Q����QD�<L�8�@�i�mhȿ��[�zjl��@q��s�~vC�8>��Fj�%V�p�BT�u��k2a�Rct�+�$�b=/��f�r�3Z� t��u�q���Fj
DK����s�����?X�Gpq�n�5vzUP�^�]�on٭�ǩ).#]�}�-E�����sՇ9���E��3,����5˺�(xŽ����M1D��1,����[EF!"=���~ݷ�u�����;6X��r���h��l���(i�p�`�t�)F����T=�W�}f�q����b���5g���_�0��YiL�1���ˀ4�/R�;5[u����5X�eI+�Ue�^M?������pG�����W��ner�@pלef3�b_��T5�!��H��l�����|��(-3���	�17~!�H�{'+@�x$¸��G�Z3H��_����R��=���C��W�=<q�'N�M�u+�8��|$~�-�HWx۵�_�Ӕt+��9*=�#�Gw��d/J��=/Bp�|��*�"�����o�2�*�`�S��3�[Yڊ�<K� ����fG3p�
P���w�O7���75t�nn<*F�N<���6�@X}��y�����{�������A��=�%��o~���b>&���IL�CY����}���97a��#��H�đ ��l\��E�����G��)��v��!p� �&ڞÄ3g��vh(f�-����b؏[Ƅ��+X�V�6��g$�H�ʩX}[0=��@.-�|���#���g��M�d�8�Nꩻ:�l��t�R���C+�����nzq>J�+D���ꮮ�}کe�:���k�*|Qh�Q)S��Ph3owi4݆�L7�<�R����g�̂V�]g���$�}&yT�@!9 A� �u�	�{����bO6�[|�<���)�$nK�a8ע7)��]|���G��n�](���K�=<�AY ׶�V{�M�>[��T�[��\�{k��ώ��/dJ�C}j�67���⃀�#ќ��>�ur�t�����*�c?��W��(��F8��U���
�uA�oV�p���/1O��-�-=��
e�Z��p��t�.
��s
��l�ܟ%H�.=��&P��xy퐋	D��ۙz�~����XHKC=���`�U��!��u���\��F.$s2g�'���0�n0�q�V���r~�8��H���=-x�׊<p�1��1�d9w�#u�L$����/I��5�S7�_�1s�EHƪٔ��(c?`��Z�q�^+�m�)����`S��g�`F!�ή�,gX� ���ݒ+'�1.�����_)s��/̚��?J	G+FI�=�z����/Q;�4��Zs`��erR�%|�y1�8=�*/��аiP�it\wH� ��G��q�F��wn)�{~d��~������x S�%`GE�y��ݪh�O�܎�J�~�`�C�r���y.�Ő$�Nq�	�ʊ岅x�ݻ�z1Z�ěC�b��/����/f�\��=aaZ*g��S՜!d?�3�<�Ytb�<c���0?���Ggvl�lE��݂C5��?�R� �@I�c�M��2%�w�����M��Ζ��5"�5�h�'ۻ,����[�|�|ϱ���|ϱ�ծ�e�}	�a)V=M8��`��Y?��9��%�6��:�*��� ��}�ب׎z��^�����cu�`1	Uk�qf�A��b#���0m�Y84lI{Õ "�v����w�N{�*[���e/��*����ʱ�k�f��*0��L*�P��C�(��=,�
�Ǧ���+�2��
��,"�� SW��;��K���Z?]�h��-]�4�e�tV��3&Uês��?>��=b�y���]϶���Ne P���:f;֘QΑ���k;X*eJ�؍��k㏱����"g��&>��n��[@���B$�4�t�E䵩�3���Y����@�]�<L;� ��r���8�x��o�2�8�c��?sP�Bp�eg�����׉�
ȁd�z�2X
�'˾��7kcpe�q���/)�#��OW�(p=�^�n�����r�#�WW��+��l�s�6t�D��%a���%�!3 �$��-�.������A�������]&�ɦ�:R�%.�˸�vK�i�蚟�m8gc/&�b��I�J/J-{��@;��\���\Y�At �:����<�w�M�������� T��H�Υ>ι�'^zF���+��s�;�lu(��Pv+f0<�R>i�4�$	O�ζ�	'C�Hj���u�W6A%��N���;��sJc��X㵞ĪpC[c��?�#2"0�����E8.oΡJ�+X�f^�#�_jլ
��. ڃp�#EuXFO�S`�_�=	��<��G��n�&��{��TL׿��%h�~{��&�� zz�+'����Y]�Z  �`$~c�����_h\l\�S�"f�sW�ąF��b/ՐOE����\��c�ٓ�g�_��K��=""��UL��"~�(��O��z9�c̹�0��Y����g ���꤉�v:5�o�8�,  ���.匆)���H����h \��i��W{��{0�I��C�5�L�a�#l�R[sG�X�]��I[(1��F���1$04�
`���Ra9�̭O�����Q$"�����(0�?T��"����XB?��wm��7]j���)��ޯQ9�5.�§�f���P&��d+)��$�OP?mvI({_��eymx��^���֡�ܲT�ֻ�շ�*�dD�&j�E���Ū����f&�;%>p8Y*0blUK�b<He(֋�-��
63p�����
0��jp5H�oŉ�Fݥ��*�a��c�I��h����Eޫ��e��������|\����d�N;q!7Vp,��qzlm"� a�>Af�o���/�)�e\������r��J���(��;�����j����L�}��W��
׌439IH�F�}�qZ�T�b�l�눿��B�6"��-�*j��t���>��p���E���V�&������*U�k"?K�8��HV��Ks�pl<i��ho����&�����4��O���K��C�{U�s�ts�,]:������{��hh��p�x1���.?s����s��vDT�ث���]���3�w`_/����{��+��=�ETMɟ���O H�>X¾O��;b � B}�&��Z�#˔�G�,���0Xբ"�48!�_�&���c�U]���=$�a ?GJ`;���q�BBHB��P��҄O䐺ض酂=�#joo<NP���^8;����p��K{L��o��w�7غ�� ��~��6p��mcW,gI�`�Ex �yQAc�{�g<�~�;��w�G�B�CG��8�Y �z�!.�`�_|RL��[��'�W��8�W��qcqƿ\4���ϲ6��"�DUqC��mh(�]�)d�z��;�mZ]���L�W/+z����g��C�C
�dm��F��Ό��3@VZ���ҫ�J9�xNM�5o�ց3���r;M�{Bc�!2Yz��d��L|����7�(�p��������ע0,8Q��?l.f��8����9y?��g	�
M`���tDN$r�XĐ¹��&O��>۹�MT��c�����bFrt�������DlۋB�^���rQӵYm�x?� �,m��!��$��*���^�OD���)UW���d�f�a���:���9z���^/�x-����\�W�Aϔ��o{���}����QC�#Á�����^�� �)�g�7�qʰ�gY���U6���=��Ça���~�̻Zx��j��<O�J��ƞY�α�B�	o4�atW;�b,�/ Br;��Pv��g�a6�`e���_�u�]�{.���J���q{qk�d�u�*�_�ſ����K����u��O��W�2�0M	��L5�3H��Q��.YAͮ*'���&�B�'��� �b!�M
�Ŏ�;Gd�\v�D�.��!U��?K�ߑA����s�� #��ŋ��\ZU���n���lLLaJʀ�N'����9#o!��D���p���jAӋ��uclp28U~�tw3l/���W����y�1�ݼ�������դS�H���چ�aA�t���Y�.oA�8���9��c0?8�S�)KC����F�Rdgd7]���.�P6��F�n���{f!��������H�n�h�{�@]�r {I�e��9Ί���u�b�he/I�(��|jO��sQ�$z�{�8�*�U'rTf�+�H�R2U�&<�0T>#���E`]?�٦�WC���[�j�(AMX9!/q|��.�@�n��V��#h��/}��3fم�/�|�N`5�����R���"���Z*7�tX��d��֤��2��&�T)���m�k2m>E�Md0���(5���<�J���;i��)O����~���/��2�6��~�O��N�~d��<��䈫��a����ҭ	�rSQ��ַ���b���"`e$X�m�����pM��ܪ���1�ʅs�b�5�2�P����� M��3n�s.�y��;x��Ł�Z��J����ޡg��ox�6ۡO�b��)XЉ�J�$w�@V5��Iқ�~�3F~B-\�z�3K{'#�Og�+��޽��������{�MF?� fh1u��cb><��g�1��3*%��!�{p'Sb�Y������j�=��3�"��:cx��Q��^=j��|OJΪ��8ޞj�D7�8��t;N{��Ҡ�l��E�3$�J���;�cL>�X5��ʚ"�k -2�tZ,A��=c�k���v�G�+�@k�Oe����3e�#��D�$��V���QK7�G�:ޙjf�}Y��8�>=�O�ёs��T�!�L0'@��촦n៣�K��w�B�
Eqa1X����6>�L)�
|��M$������Уż��b&?�t���U	2�r#�0�DW��U&VtVk#�5��Ui����a�STѵ��[ւa�4�3�[�@��r��D�4����K06�@�礜��ǌ�����;YT�2I,3��̩��Ō�'P�����*o�ķ�Y�`�KPP6���8�E���1]����d?7�A�1������z�;�z��ZN4W�CZC�=ȭ�:Nn�z�Y�U�w�U�f0��.�����%Y�u�I��j��`R�7�ѪOZ�s4��
D]8�8x�IW)p�?`
�]��LU�>��"d˗g���B� ������KH��4x,��ð��$㤩&��[�Q8�|�R�{%�[g4a�	w�]1�[�Hh?��Y�P�<��2Sn���I����l� 5��:�0*ǎo��H��/�2�r���� ;p_(x�4R�h��QL�E��n�����y����z�
|`!��ǃ��m�y��CKJV��rpP{��;_�q�61��@e�#fֻZ�6���/�[x�D.a�QB1�-���Y3�d]a}
��p��BKEv��ˎi(��dJd*Q?��՘ə�GJ�ґ���r�%8&�TW3O���T�M���/��%����Q�s�h9�/��A�OW̌s��O�F�Ο8	"`��Zƴ��n��fܬ�!��+�ந�UJA��RpQH�����?>��GPv�͘+U64֡D��nFnp+�s|�1�Aڧ�d���G�<��d�^����L�l�U��|T|S�����RE9��Қ��5�V�7˼:Ýrq2g]cZ]4�AJ�~�������`K��޸�o�if��J�ظ;�w���^
��eg����*\�ԏu*�%��� H��̨�t����7e�����0���%�Q:� �E/��m����J�+�N!���G�<�hw�|���� g�Ƽ)ö��KrWlS�=���~z��p�T"�j������Ŕ�q�~f��(� �ם���;���&�]x�����"��r�$�2�=�o�Y�._dG�ʆp]�f*,Z[�Z-Lj�����O�@�[�jG[��yR��^���eb�_��(&*�EA]̽FqZ�����췊����>��VT��^ U*h!Mh���Ji2!iA6--��wJ4�Q��ͦ�G��bu��7+:��q���k���*ԯ��!J+�~�t��xPy��a�-�����`� xٸ�%P� $=�BE�)�7�x+�;�@Ig\Țc[݊��.x�9�cm�q�,+\�������ac��Ǌ��٩�a��B�l�̭;MiH�Q���)�cş����G�ɧ-];�d3+�tgTt~�)�gBǉ��5g�6[\.��@҉
J�l���E��(�zZlK87ƌ����s�4/��]��������d��&�����۸���&��Fo��(�\����/�J� xx�Ç-�E�mm���τ"�`;YQ�9��H�k]��INE*w�4����9C�e�W[)���`|�K�T�`����n^n�\�?s���]�_��5�rtdQ�(��Ɓ%UK��d�,Vb���� ���.��Ms#�������7L9�B��b��3�����S��j$�Յ6�����M'��v�3x���!��7f�3<m
���=��B�pm�h�� �ٷ�He	*;K�6�YKwj�uiz�*M�{�U>SX�Ah�[$�*U~��3���?K\30��`�W dϷpih}��t������;�w��5e7�����6�T�[ޥu�p��o!�?å��
��
m;�)���7���3x�0O%Wq����_v�dkId�\)�C��'��]��5��!Y�~GG�����baa��WF��{�M��n1��`]�TI��&܌���y���i�opt�F�m X����k���n;-ǭo��=���k�����)���,���aD�0蠞멥��%�o�r|* �Hl��v(����;����sQ���1B�	������	�f
&�9��i���EUD�|�(EN��=�(4#_�6��Q���m`�4�ah��=��f~����=r��4�l���8(�������q�`u����5�NPGW"���סq�Vl,y���,/(�������-�d�-BD�ۺ��
��6�-;팇�A(?���-�:����O1OF���k�O�d��X�"z�9� �>~�q��PEP��s�;�C��.f^;�X��p|
����b
��:�H�`<�%�������S̉W�c�f1����7�Ȅ�E&:]�t��kRv���彋��@���|��YN� ���Y����A�D���H#��I6Y���ޏ��p��\GC`���Ah���������淚���\_������Fj��=v�&�2��wA1��L� �~�/�p��T��/��iS�^Q{�L
s�7DŹ6α[a��#�j(N�B��27��(�Mp�G ������H�S.��pi޹^�*?��A����a�L>�x��9_ɲ��#W;:�������%/6Ʈ�x���C����O3߫_o�O}��bFOb��_���$|X�������-�(cp�}S�Ls ������
 U��)g�;�K��*BZ��<�˱��+�#�(8y12�cK`�6�~rd�v(�s*�,ﮞ�n�����|/��"6Drw��f�#�?1.gx�L2-�LB]���+]x2��as���(����xJPA���8��{P����Щm{��a���*� ���a�B}ɧ *�*��H��Kȝݍ�.�9�
@��5%b�x����O�|S[��D���KDKc)��-KP��頵7�/�����D�{�a�9�p�P{1��~ɪ%������^��K�yһk�������(<g����)��z0�xy���4�0�g	E����,~�`�el����r�#������k���1��uǔ.v�p}|N�<�'W�s�Br2��3�YB�T�ے�/�M��g�'Y����b�m�Ϥ�����H|B	�?�\�([As�Uw_ѯ�K�8�u �t��& ����|�t1���Ӛ���VZfgb���Y�0����j��^7�3�r�_����Pz�|���Q��U]���s}���&0�8W������Č��H�L�C��>e��`{La�3����X�j!���|r�G�/�h2���� ���L�P�q>�3Μ�������j'���]*0!H
�����@4&�R�V�D��)�W�yƐRf����ms�M#��1	�=SX��?R�dE@~>/$�g��ҿ�+�r]��KMދ���ȇϕ��:��|�1ԉ��2_�.�F��W�Ҡ�����Cb�D�b�}w&�@���oM�g��6�+֤~܏�C��=Ƒ�����(^�ae�X/e�\�~��%��`�}$β�% !���j�ΡM�5,���JH�
 '��-��[��xb�|C�S��
A�yEY�?�K��l�)k/Mۻ"�O��!k_�T�����6�L�M>�T���# ���q���p)Ps�[z�ǋ*��a�.Xv�䘱<��PG�>Q�3P��r���;��֛'kQ�o �j1�/�O|�d)y�)H0��?��B�ih3��2	��$�'/9�B���p��\�}N���4��1�����:#�w�a�9�y����-�V���ިA����Y�5�3��c P������>����c߂:W>�Z:�r1+�3	k�^ԩQ��fɍ���-V�\��5�p�_�h��eE'���#:�Qj��JV�~Uhn��ܕ�����'�#��+>�S4G5�HSZ]�3���#gW�+�5�e�D�#͎@3@z6��h׎�-�uSc����dC`�9�oƎ�p�XY��ll�}XF,��M��}����	2jƺ�WA�	���>���WʣN�な�['p�R>.XnM���� ����C����S�|ss��$���т���e�`^m�3i�u�� �߬���5/`S��i^i�?��������>ω�V���H�*���d���яc%�b{�� �����7�E�Nac��r�1j}'vtI@��&B�a�9��U�PgqR��jd�����A�}{�iKRm+q��x
�+���{��%��_Y���s(��(�$YD�?�J��S]�W�-��u�>��>D)���Qf�����ύ��CĪ-J��+��� �I�ݡ��~N�9=沩���x��b�r�B��\�qg�?pA�L�	S��.����Z-�c��EkB`G�e����&k��ϳ��p��;BcZT������;�����Vv�`�bp�E��j*f��>��ʖN-�x�%�]K��'��;.5ϱs��=7�٩}`�z�Z�5��?�α��b�cf/2|h�r����)~m��U�w!����_Z���׀]�QW�lcNE�עH�����-�G�vԌsg�ڰ&��e"~������h-(�W�� ����ܞ0�_�CKW�޻�|>��+ٿ������K�e!��B�yU5Y�[!�A��.��>\���GB�3XU�f����]��@��G'���4l�8}�'3Kz��DP>��~g#5���b1�@� �|Ţ%��<����7���3\�pld��:[^�ME�'�iH� �<�i6\�쿹��̸�$�1td����Jc'����ُ�D��=��"r�K����4�]H]���K�tO����\#u�b�L��Py������%#h���L.ͪ��	1�ّ���t���j��7[�R4�F��W��,j��s^��yhK�*�{S��(|�V�����-���o��;�W�7�b匆D[��8��h6؀}�F�I�qU� ���U~x,J8Ä]��_���L�:��NG�����XD!��6.�]i�,��ف�|��:[���L7�Q���`m̉kA�����Hz�?��@���Er�^0���W���4�<R#�x鬃����F�JC��lCE��o����pҙ2� <`Y�99hU�e�\F�BmN<��F�g�jçi��hk�R�~yr�>��?�L6�`&줠����M����-p�1�D����vO����;#���
դY@M�`�T� 6�1�$�"u{vd��n9$�/�)=jT_D�u����(�`���cO=%��9��eԙ�$�!�Nf>��&Ghe�x��Nh��ј<F�۸�>���Z� K��sIT��*��Ҭ��B\":4WK�+:���W�;�����m�%���-uNH�(a|jb���yiFp&�L�̶9�ć�v&е�D;[�K
����uR��ț��W�Ô��� �\���w 2u�[�Kh|O��]�BZ�-W��X�m��r��Nli^�?��-p���n�s_s6���0�M��,���m,���B����hhXLu�Kݚ� $�o�p���|��5�N�r�jRd9wn��`��<��)�o=H��Y�F�	(oQ��\Z ��s�Ş�����;�`�"c�[�*�{GopZ����p�?%�e`s�蹜 �ƪ4�b�ʠ��k��eg����CZ�Cm&e�G��^��
K�=1)�IN�73NO&
W!1�ñ8��)2"
L���r�VM.f�(k��|�|���ܤ����YȤ��Đ���Z�ȟ0�I�J��u���a$dY�-L!��+��Z�_�vxk�n����Ŋ 
S˜.6�W�6ci�T唍�k�/�Q���H������N���ӏaT����y��}Oh�]kvTpñ\��䋍��B��D>����O��3�Y:N�2'>�ky�ġ�dc�N�h�_t�bgwDV��\��}����l:����!��`3@n�o@��=�=XѼ�y����.��z�@������$;��x7����޴��{�'ю���qĪ��.�8֓�S����̙I���/M?#%��̻e����z�X�Bg��J#7H����h��
�@�~��A��o�@��;����_�6s���
�bn=W�(���d��ߋ	'�Ȋ��)�H�����G&�;�AU��2`A���b�yO�$�t�Ρ�ҡyy�
�1�
�+t�e�E.���i��3~��~�������!g�J���֋Z�8=Ȋ���mG�2��o�KI��Jf�Z��nD�W�JdKċQ�
�u�Q�t��o�ܟN��5�2Gl%�ɊB�q�ށ}^,#�P��h� ����`��?8C�r*�Ʋ뙺57�}r��w�2w�Dc4�W����?���U_+� �F�\]�X���E�i{����.FʨmDIL�J��`uM@a	�aH��������f���� U����%%�ȖA������K��2��`e��v.��,+�U�8�f���:}*�*f��MNWxJ�
B�:]�NW|�-h������칺���,�l�X2H�i��S�J)B�`�ղ�[���X�	�M�zc|MUR�F����$V���� _��3dmxS,r�R10{'eZ�¹L3�?�yUl+��ȣ'���3.�����-ƾ�S�Ͽ�S�-�z���JO9�m�g�m�T�� �]�3�"�܌�e�Gm�R�Zd#+��L��Γ	������M]�R_�H���M|���Ł2b1��A��H��%���×�4c�t#�׭܇����*��)�GZ����L���5��ծ� <*�/0�Ԑ;}@)��Kv���C}�{�K:�Lpv�SN!"@�٩G/md�n�S��*y��6VW1�j0�uRz�yb�f��W�+cf���9��=�L���g��@?I3��8�A�"Qn�'���HĖ�O��)`��eI��4D�VGmZ�54��zQ�F�U����nR��Mn+hf7������n&�m^z�P��Ύ]M��O�[��v�����S
�7hl��Ww*s��Oh�'�.ُNz�.a���>P?�g�LΥ�G�(��6�cׄ�>pŖ1z��f�xr.�Hӄ4�֩���w�]�hc���l�s��˧� �3�w�%����0�O��w�̒Cu�R+C�T
�l؟8��L�32F�y�s�&)�7�kܡ�-ۥJ����&޻��v�D�^;M�A�=��dp������.N%U�-�F�f]w� ���;>�r���N�)�,<Xx��>�n�e2l�+W��,�X��]�f�����V�l�3WZ�mA�;���R��B�f�s���+��u�O�q3�Oy����a�{W�ě��0)?|�+���U��M��K��D �V�$Q�\�i"�^ݫ�JX��7�pi�:Rd$��w´��;���̕���:�sӆ9�b�p�"�~���5�U�Jn�}O3RGN�xK�{�vU�G���A0�]<�L}�ݲ�P
�?oc��\M���hC`�*/0Q�����-�\��a<<s	K� -v�����J�7ю8>_w�a���{�'y�����XYr��[;�d�[�C���\������V������{-[��z#���}	��p���mw� 9|���a��J]��R#�8s@�@0�,m�d(e��M_�����$E�R�U��`�8�y,��-$�~�{���:��r/*�2��#lY�"S�L1�wf�Hyu_���;��Q(�1��t�e�?�ٳ'l'��н?���Q-���H����.4�����=���+�����hX���oL՚����)M����ֱ�s���V�r����Zх{�����1�'��	�k��4�+�TJi�J�(��S��X��\<�����Qp�_e� 0[�ì/i �����O�����E �np#qt�G9��#L���l�MՍ)&~��N=�@E��0��|.RqD������W�.iR��2�}��R9�?�0s�l\��2��|m�U*hd�x��U?�!AnZ��4�#����`�C�D�K�j�d�o��
J��Gc��q���v"�5�A��3�psw	@��pvwL~���fO���}�T7�K�E[��=Mw�����),�;��T����g�h~Aa����߅��I!o^�Z�_�@X4���5�5��Ϳ0I�Ir�����3݊�Ƚ5q��'r�Hw�}��
d�Wi�*֎��{����<j���8����>U��� �0Xz��d�����y�ѝ����k���]����/E��1��EK�Z7搖G�!�?Z*-zt�T�$�P����H��H�[�A��x��na�5n�TG��)�R��,`���f�� �Z"ړ�<η6��vÀ����'���\ѷ�EJd�����L��mc�j�p�
�Zozl��Z��
��p��<~j5��Q��l7�3���xټ%z���a�9�(�s��ϺBi�/,�������w)���G�p�ܡ�*ԑ�a������~����V�jiI�n4.`�E��w�e�J�n���p����~7x�^�-�����`��Ҭs�y���܅{e#�Q���h	F1�ao�}����g�%[���`��h�K"5����oi@�Y��Χ	�o,7�V��N){(n%w�ǜ"W��j�Ŏ@��և�u{�S>^��A��1D2K[���Ll�8_��שi1m��^� mK��vFT1���������
�on"gp\ ���ܝ.�����>�Ds6TŠ�P�-	�s�	C�o��x`���M������[��+��;'t܋�X�ǣ�A���K������]���v��J�OPͻ;��������k8��n��uUi�?

��2��T�t���'�0��u��'�~�L�U�����g��b����M�߽�v~��9q��jr5E����S��rWL1T�`��x@U�6���G���{��?�$�@�^�_x�<@/�;��6YFU�4̌�/����|�����+��M����I�ӭz��v��:��8/�&ɐ�ʥm���)~����C��H���RP�����v\ݘ�2�~.Pf<����:���^�EB*b�7f���eoxs�v�H�`�ւ�ʡ�;<k���ٱ���� ���W&��^E672 ���+��Q'��G�?N��P�����`�&9�I5�Z+t�1�dB��/���k���3����Ŏ�Yn�����;���V�l���0j���f$��S�/��3�[҂!Y���^#N�-�k�h�k8(�׮|U��&-��RF��V�d��d�p�(&8��	a�Z&ޅ�9EB�.��y��XUr�+�\h,��k������(��=}A��U��M2�_�f]U�*� �bO�kH"�J������l����n����n����QpN�jZ���BmӉ`g�(a~J��m����	��~[c��Z�g�ClK�%H�4H�J�;Ɔ%�bP���4ܖ��F��Uֶs��[Hm�l���B�Oh�tPo�x��$#P:�˼�X� ^F�~�DƩ2-op�au�� rZ��gl<�M� I�,,t9�|\<#��m9�����-����Opx�G�a�Q�+Jh�a���U��~������2����髳yҍ �"#)Ʊ�&�&Һ�%���r���5r:y�t� 2]0�A^�k��:/�[r���ѷk�q�öy �$���Ag�3c�`c��Sߵ����(�ZD�R�PP�+��S�o�x�E6�������lz�7^�l~���v<@�����3�@�%���+�=��6e��X�[9`N�1.���N��k��.��� �/%�ՠ�UAI�t��!�Us[o�u+�Њ�@�X���D��e�f�5yG�]螏��M�yj��09��Cn�UP�3�5S^t�W�K��i���P��<?�M8-�Q4�r>ѵ��Y�^'��~�-�jk�@/s�� Z��.X��a�����,n@�����ުk��)@S`Yl}.x�_Rlɱ+��ҕT5��Ef��B庾ۛV�X�����F=yJM�q�������,�V����Y(o�0�.�1y��bs�0��6&�캶t���/ ?L�����mu<��Y�\�����Q�{s:�	f�[cۄ�<�K!@�pá�͓�l�����B�K��%����	����B��x��I�z&����!��.�}�1���@�0����� �F�˩���������rZFF��J{k�䷶Tܒ�ho^yk߃�'i���KHV⮭�����>�������v�)�h��)����x�˰G9�r����zA+��H�[u"�4���kmȤŖ�a�7\7��'�N*��/3Y�PCS��)0��k�͖���J>��D����%Qi
G��aK�&/����=ea4F�>��%����`�0}31���m��Z�*éSAXų�7�cH�R{0�Z���a�=h���e���Rbz�dk~6��!�\��~ϳ�{>��􍟡��˦�a�k�%��#$5��s1z�s~+f��m��`а�K��Cl���>D����S�}5*:ކ����?����+2�����4�t�].�nS��o�]�l*
���,��獉��n�W�������֥��ף����܉X�2�g���ק/��Q�ﶰ���S�xp{�Oyi䖘�K?���5����J�!���p�]l�T�)�~fL��Y7#�ڱU���/�.G�b���0�9d�$�e��4��3�� ��<��� ���o)���G��Wߊߡ�
 �*ϔPN���n-��󐷃nd;h�W��@ih̆({�a[2�񏌬05���#V�2�-����q��cM��AU\�A+P�~���� ����cz�Ui���wv/��\��7�l�72���Z�E�Y�\��,�6�����9N����"�7Z�%�?����nV�:3N��P�)&q�{�e*h*����F*y|���Y^E���ΰ�&HE�|~s�T�}g�K8�r��<(��k����7���_�l|uE��8z^1!��°�y�l�^T8Wwy(ZC+^�c����V6[]����kH!I�i�v��%Fs�?���9���l�Ϯ�GK�dCN���h^b�Ғ���~��c痹��= xb����I%߯d����:U5-�ES-�H�!'U�ֶ��\P����� �pܸ�YoBt����t��	�.���>���^����Q����N7��Z�iay��^�z�'9�4�@k��u;�x���ۤ
��:<�Kb�-��_kY�Q3��i�6���`)|T��*.�P�E�x��g�GC��ڕj�N^[>h��ɧ�������'2,M�E�f2�[G�t��� d�5�"�%q�n��VO?e�~����ߑم0�@}Q�c<���k��3��w΅��?��n'��x��}��v�[0������*��</�5Edvעx_�z�\]-�ii3&¡�\�p��Am��{(b�v�7 �J���D����`7��e�`�� Έ5�ݱf��{����������dS�cV�������j�;L�ҒP��/��P�l8dՎJ
�q�Y&[�$옜ou� b��
��u�4|�B<{�$��ۀ�8���]�=�4��܏��F$0��+�G�_cr�Z}sUI��o�8�L�'̞�J�pa�q����ʝ]��$/��n�x���"n���a��K��l�� �a.�
C��;�^�܉
��Y�y�Y9qw"��Y����޹-Sv�T]�u�F>��a[s;��lA�ȏ\@?+�R�\O�����+��J��v��GC�2��s'/��v�h�� �W#<R��w�,�+w�V�gH�aE&�	���"1�b@a�\��:����5�/��5�`\M>��ۻ>AD��b�7l��!=��"���_Zǈ~���� UV�q���1;iL0����5]�Y��&�6����J$:��{@�lc؛�H�j�E�n����
����x���������0�&�<��|�)��jS���ڗ��0�?�[�#�q(��Nٔz�@̀Ӫ���߼���73'{l3���Ŭ!��%f%��t��OnA���HU����'m�s����,w��~Ȍ��)<��zU��i4C��'����k� ���	NrƏ9����`�N�wA��iP�R:Hl�.�h�{�"A��K�im��6�v�� ��,6�9�q��N�$n�M����`^V�xw"�-��"�|�A�?>D���y碪����q�E��m�i�L��wBVr{�72i�[�Cs�:	���$W$S�>͖T 1xZ+(���d��ln�ٰ�����{�׳��wU����<��&��S\jH8ܖ��e��r��x�V{�����HF��ُ�|*��μ�42wS
S��������-~L����������3�S�gŉ�Y8�o���>V���,*�v� K,��L;���P��j��A%�8
*�=]������H��9�_n��m�8gȕO���A�l�<2!J_"��t&�u[��ѕz���)�p�c+!�V�}6������,������)��ݩ��v7�E�:Ç<��-�mˡթJ��b��5�Z�4=7�k$; �36[�l7֭�'��,�S�5�H�x��mܗU�p�ƭ�����Ap�'�.H�q�/۟�!G�EMJe	�S�t�� �l �	��A�[�vk�b>\q��Q��J��p��E�����s�_m!H��zoG�n�kN-Sx1�)N�Yq��h��Y��\B�Ѐ����hR�Ϸ��q4J����Kê�T��Lc�����#�h�D������������:��V���jzN��I�a���i����G���j��T�ԩF%ɷk2p��Ks��ɟ�ab�1[�`=��U��]��w6Q�ꆛ���p�y�p����=0�B���
�X��%\�y0�Y�dh#5����mM���&bȂ,4�b0.�H	e6�D'o��^���yxj�Z�>0�	��a�5�Bθ�z�N`�a��Y�h?�O,�ЬKwC�]�OS���^�/�Z�\Ǩr��t9R��ǫ��o���J�E�-�����~���_�hi`i�	ZW��G_ݍK rtI�06-����@Y��6����J�,5s2L�6I[H��{��[/y��2:���d�.G>[�%Y���i���ѽ3G�=Xڴ�)g�ɑvE٢��	��CT��5**�O���oSS��"�f�tH�+�Nƙ0	�A#�y�@6����Q�q@E��Ӱ��5�{Q�|����BgJn͜T~6�u�A?��װ}�-q,��$��Y�6��9���e�>�2d�j��l[����
6��y�R�*�����TMw��P�r���������3U�}7z���=.*=��z �|��a�KG��(וpD;��C��Ȃ�՜3e��IB�3."����X�4��艮���'�@�" <�G���n3p�@���u�l6���3���ө�l�9 Y����-o�n#�� �bBC5����D�����)��x}DK̉�W�}QU�l�a
e�>Wx���};3�<=�=
 L��q���V��]1z�Ί�YzTݡ0H
)�1.��5q�%G������Işt3������ص���dW��+)T�e�n��A��44�\C�TR��"��;�ژ��<����R#�U��0b����q�Na �X!���R�
�FFxh��`�/4����8Ռ;)e��q�)�_���� rka��(�~�q�?4mԨ�r|��=�z�ê��(ά��՘Ĩ���D���y_ٶ���e��㳉Ui��M2���B�1�����z0�y��c�L��M�G�$]�6�|����JZ�������g���y�9d\zcJX�YmU�XW6�c3�z�م֟8�,Y.:P���_[`��d�����#�)��N��Z�����j=�����
�fE_�vr2���Nq#QR�j`0f�I���ۛQ�D~���Y- �D�6�9 ���$܋�k�I�����\\>K��饲˝N�I3�����{�t����"�����W�kd�f�~.&n0�gl_��v�֌��$h6f�}�@��\`�F�A��|�ҫ�[&A��� jU��sU�r�Q�-�s���{w�!�����>�G��e iw��BM`�	vN:.F��$_jJW9O4�!ݑ���2+:f)1�D����0���{�i["���t�@�����N��BJ2M&�^���ml�+�\��׼�x�C]�G�	y>~��W�/����6�����W ��W9��CN+7�Q��8��F��/Ъ�}w-ѻ85��~�Q��f�-��~���e���bE������>�t3u��J�`Z����
�ޜw�iS���]���`�+a�I{�������fE�k�Y_���P$��6���*.h'5!	oĵ����Zy΍f����s`���YS���� Z`�'���Ġ�a�<E���=�k%��ɻ%V��^E�L�\�'B�!���Q�G����x����a�9c�0�EC�䒐ǅ1�I*Yk�H�h��M���N���N��E�rJVZ�;*�!�jǂC�q�ΤZb���ִ���Y5�Ⲱd��F�8�b�Xh�+������P�J�s��e��V�R�P�ҥ�,�a2kF�o�t���H;R���b�{���w��k���ݜ���_ϳ�:Q����Pu6�Om\��>u�8�i��x���"�Q!mħ�t%�&����)H}���;����:��9}Ҁζ]=�ҫ/�i7ŝ�H�?����Jo���ōI?-��RfS#�Ǎ��^��S��&,I�6����d?��|���c9�q�!~��F�pS)UW3^2f�!"�<��;�ܚ�5��V����_&�>^��'?����G�+��}WA������������YO�CQ�$�����3_��zǞnT :���: >B�Z�{����f���[Rv�j���յ��#�C��k�l���S�\�b�q��V�>�6����z��D3�%���BS��K�K^��!���OɁ��� D���r�ʣ�&��Ì�%8�4 #]�sV��}�O� �8e^�_��H�T��Y5�4"����F-u�lV�7ʩ�e(O0���J|��q�v��6��)�ժ ����h�r�l
��Z! .R�k���-���Zِ_O���z�5&E�).�d�+M�e(j�"��{7u�� ��9��*ٷt��{���I��Z@����	$�v����\R��+y�l�y>1�L�����퉚����{���n:%�|I�`�8&pU��|�Ee�X���n0�҆�ջ���26�Th�x^Dq���ߊz��WS �"����:�X��磈�=?�/�;��`�$�g�8����?,�K�`��w���P����a���Kb����Vz�v���Z*���I��-�x��Y�%��j��N��������E��
 �����!���it_����O�M��v�)�9�8�6ɗ6\�q\y�'i9-�U�6�����!�c�1�>LL)���㩀���A,��s��N��AI�+Q�A��f�rT=�#�<�����z���J/L��ի�+2H���/�"E�ޒ#��W?S��_S�K���"��p��/� u+�@i
r�o)1�~���D��W�d�q�E���3��|w-GhOJ��*o���Tӻ�e��M��K�|��/������Q&�J����+9�T�3�<#�EQ�d�B5�^�9��R�v4)fr��bc���eA�E`.K��;L!ii��u_+����:�FT��Y2"��@<1<]Z��������0s
�t`��à��I�.�[��m�	�Q�掶�3���]%Z�ٸ��Kǵ�ٔKH�n�	7�IGw���m�8F�u���A����f�x7	�1�|.*�L�w>�M ���?_H���	��d�ﲬ�������[a{�xyb�&��{��6��������T��D��]<�<�J��ͤ�C_2��Ӆ�˝��3�WoԖٝZ�~��9�����}Ij?d�GUo������1�D����������@@�b��h��u&�/8�Q�+�3O�j��V�*x�O}~����S�F��gAZ��0}�Z`���ܠ����E���9�&�s5ߣZ{����@�HH�9'����էu�g�mXF�k��yƧ�����݁z��M�!.,��71���F3q�턎R�������8��3)��B����A�N6/<��y����sQ�g!����I�OkL�ٙ*:E��&��*?��m4D8J�t��H�o�FECJ��)aBt��ZG�r��o��m�#���	��!ݘ�.�
oAY�q}��cK����Tm�������������ZX�`ch��K�R��+v֠bK�4��`G�R�@��/ǿ���{$�'B�����>�_�4kv?�x��E0'�4b��~�HM<�w�J�@���!8��W
��&���
�<O�o�� +�'1������WB�e�o��ߥbŃ��̅p�'��O<�{��lC݃=�T/d4���v�kzܵ�[�r����#���,����������ծ����*��z���6w~����s�*=IL Q%K:9@Ĝ�f��U�fX�٦
rw4sv�VnR	�ĝ�3��E9zk�3�u��mg�*��0��K�[^���]{!�����5�������N��u�����$���U���V3�M� q���bK�ǾPqI]'����2خ�5��9ʮ����4+��?�� e y*��/{ږ���=S.H��0�@砥:�. ��#@1"J)muD�/���~�
7�}�Y"�r�I݄�ݐ�w
p�}��o���ۣ2��c6M���O䰗�W.{�)�WQLtu��ʘ^~u�(���,�.�@�=�nM�3��!�M�G��}��L˺�\JK�o��ݕ�� ��I��8l=�U���9�:�U��qu�䌑7���(;�v���(���2X/���ʎ�i��K�R����Î��\q����S�.PLp�i���z��*�����R{����9A�:z67�A�����+ˈ�����N^>`\JN-U�/�ϊ<Yf̪�x�0}TE�3��`+F�N}З1S�LQz��������#⡧b�Vhg�|dDdS�����$���Lf���%�td�I���0'����q�$C�LQ?�{I�l(����5]I�S y��bGψ���׸��_�]¢!N�q�U����ȝ0�꩹�I�����h7O��K_��a>.�k52S7\9��W%Q��$+�&Ħ��D��ht�u^���e`DJ9�U���c�})�`M������ʿ�ʂ� �8���݃�Ǡ�P��j���2aq�gZ0iR��ŋ
�A�٪
��beZG������.?%;�4�*�W����m��jTu��|$��`U�}[�i���,����_��(>KB��P"����
耘�?�3��g~�T�0EA��ՠ�s���m`8>q:���Ċs2��;W���mM�g��2@kSKA.m%���_e1�����ƽ��9M�{-��4�={��H�����!d)JObg�����E��AUP����)"�tX���)1B��1�V�D��U�������_���@�����`mv��>W�v��w�U��MztD���p��A5(>~��_����`L)�����):�~N�E���;J���ly�L�ɝp�WN~���ip� V9���z�Q�q
 �A�9���@d������xPi�V=�+ �H�B�/���g Ig)h-�W�Kv����3X9r6>�X�mrv�x�4�'�7���5� D�4Ap���&)��۵���*����Q���m1�l}H���W"V�uV5-V
!m+^$D&F|�z2H�g�0�/���C���X����� �WL{����/���}	dN���p�?ӦG�xiL�ga�,��m}7��]@e�b��](�?���G�ix��0���9����k�g	����;Ǿ��3��h/U� vb�^r���n����}��!l��}@����*��[�C?ĳ�Jr)�Qej�^s��h̰f�Y,S^,�a �~�-U�_D��$�X�b�Tw����*.1�M���r��=��Z3��^ >O;��U,p�v״�$Ρ�Lz��f O�Z3Fz�I�w!3&?]� �m^f7��U��BO�b�U׆O�M�(���0Օ#�%ܛ��ϐԾ�TH�������[Z��3Q$J��27=�v�`��
Ti�RJ˘A��Zl����r��Ԥ�;Ny��u�&��6���O)[�Z݅� Q%�� t\�ꥻ����h���O���:�g�:�Umn��wHd?�;L����Ԡ%��v|~�=�fؾ��6�@��u�q�_�r����sN�f��`��:u<�V͇�	�%���]��lڊ�I�A*�$��l�-DD���^9���6��[5���M��j5s�#KU|y+O���ըDR>��ղOH<{�����
�a�V���
?��"M(I/˅���v�W����6�����P��ڕL��|B�x�=$wx���C��͔�
M��ܽ�篸��`����{ɽ�އ�484i��|���'	�
	״N`e�������֍�R�۵8[]fo�ĵ!�nG�v�P��C?o��������?��II1ACNL���p\6�aB�D��&��Ě2�F���Q�"1�_X���>ez7����Qe�v�`A,���V���d�m^[W(�4(k_>r.�!���5��]�{���w��ތ���u$w�E�"���z��1� 3a5ɟ���lMf'�m&����Ty�b�} V�D����ׂ�|k��F�2�4�U�3���k�?P�h#MOU^���.=�W��R���7�
�J�^��ؼWQ�]!}���@��V�Eh~��?�B���ܳ���y�E	J�#*7x�����S[`�d9Ļ��H�Z��H̊����n���D����,_��x�g��L������9��o_w �j��:3v���C��U�ά�m�P���Kb����\^A�r�إP?��>�����9�7 �L{
Dt�=\t v8ӊx���������S�bГxh}|��!��M���ю~�W<x�^t&�H`��}?�>�V�)�:'MO|;l�aA�Wls�e_�
%G�y� Z���u5��Z��ޣ@�x����Q�"�N�_Db�x;jq��p�R���d�t�ey+]%��5S(�Z�0R�8�B �]�N����M����e�lUQ�w�eg����,e�Ɠ��Gn��Y��5bP%B���q0Sa)�i���Cr���h��nP�M�RCv�Ӫ�Ky��y4Bٟa�gG\�=M"�I�Im��!_��JQ��!;t�s�H-�c�v��'�i�L�5����|�}�ht�5j�#�w�*��XQ+�<tLK߶���z��H���d�_45�.'؄�XTf�=r���^��H��Yo�S�6"7E��Pvbh�������*��Lݡ�)#�Ѹٱ�b-?�f6�5�1�a�~}uJ��a�ϔ��b��j�{�|E�T)�S����t�as���O0�n�X�j3�^�T�ow��_sOV\�����"นEm�H��A鴡��@�:[�N��yסe�a�ؘ�v|Fu%h[ãFp|�j�H�)�|Z���R}��.�B#�'Y��2߀�$��bC���V������PT�D�#�	o�V�������$��62�硛Yw�)}�]��E(�]F�'L�i�@ZA�����N����i	�C�q��J�PID.zi����p���%&!mB�VJ�(����)'$�e@��\�lP��5
?�3���I�T�sM�N���K�O���²X��-i~=�-1����h�R�L�y��e��q��z��Am$���i����������u��ڬŢ�޿�$�MB�s��@�ە)��"�Q��x������ޚ�i�+��o4�ݲ�ZQb���7nP�~����zD�=�Y�3<�'���ZLu�D$�E�Ҧ۵�F�=�W>����?��9ώ���ER��=~!DV�����EƷ���D�EB��Fy�&��������b���(�N[�K�Dr*`-_d2M5��
�w�ōE��.���O��2��&��΄���v�������G��U�S��l�IE�)~�jt3;.y�[��`�W����CN֝~�H�*[������D��Kz��W:(����z�tG�JH�IT�u��\$>�i*�A��Uھ���G��6?:H�����)ŭ�Ҍ���~CR �P����ƽm�@���!���8�����,�u��g=�oh����H�6~;Y�6Q$go.qs }N��=�zW�(|��W�P��N��L�H���/04Ȓ�F£��{��ҙFӭ�Ӄ$'�ʊ;A���Z�w�����z/ȩ���D��eG���~�sb�pƾV��薬Ζq�������7b���eI��@_��������a���}a#���ے���ύf�c+2�O�I�^H)ж*�x��W�����oz+��k��T^�3ӕ�'�����	J�C�� k���^n��!K8ʚ���/"����tO"���f��儎*�^+�&��D^���!G�˾�o	�H�̃���p��m��̬ݩQ^�!0p��/MVJ�r��"�C�>�����m9db9�5x�dJK��j�s�aQ�ix�2����+� 0�%�	��v$��̜dW���u�͡R�[�M	�U:f*�����g���XIG�\'wY,e�����"�@���	:X��~��a�������FJk̗�Ia_}>SDw�L" �͸��J�ޯ���Kk��M�=92��w˨��D����ݨӐ��R��\���-�����,y$���e�ʞ�؍41�R"?$�h�� 
�"{D՗cmץ(mte�]|c.���`#�L�}���2ʉ$�~�� K�|O��,�#���˚���&�����Z�D�Yx�������]�&P�5j��Y5�Z��?��`#H�%��+�twQ��Fy���z�x��/�V6��Bp�h@sHE8��ؔ!��\�ҕ���7�6x���ؒ����;{^X��QI�U(��t=s�������]ϐKvQ�f�������͆(ա�})�H������`��������B�]F�tL+r��f�k~�ם�RxsI���� �x�����c�T�"!�{���+��� ��y�4E��m�j�;�����g���q���1f����mȈՂ�5Д�hz�]ylӰ���X���84y#�6�gK�#��?1�u�����7-��
�i5�r[I����0�+nۺ�ל�^���9�i�*9�S D����\�h���ш�Q��JQQ4N����m%˹3rˏ�����-�|��Jl _BċC'�]=�]%gKG�
�;G&� a������8����Xek5�� �Zz.�xm�ip����6q��Y�E���!�)�奙3�Āx�%7JZ��
�z��vвWgd�Y�������=��c W��_p?��;c-2�F���g�i��%�*p%v���淽���)(OY���>��K�	^d�]	Bs�|d��1t��JO�W)k�>�DgM���n9�'�&�P@N�h�0������u���3y�F.��2 ]�N�O�`Ҋ!~��X�a�PNU�Y�nB�;+� -w���t�5-�W���'CmUK���F'؝���f�Sg��USy���S���*>L:�>,�ܦSSpF��KN].���Z S��X��\�;әX�캡׹�U�B�7b��\>�g�PCX:�Iِ0z�1�6kB�G�Ѿ�a��d�o_�.;S�����έs���d�VO〷�«,��kbkX���re�Y!M�If%�=J��Etee�S ��w�[�)���� �ꖆ�z��	����`_�`�JQ�+M@����Zk[�ܩ���kD7P	�}*�Ě�{>3n����oHs�ݩ��"�l��#� �� �rmM���J���R M�H��~P+O$^�	S\Wjs ŵ~�k(�$tiN
�1&h햘�u�A�lѰ��l��u?zs���*���JO�>M7��d��qܴ�^�r�泚�.0�圚^���A��2�D�g#���QI�E�!���H�Qe��
�*ka�=�r��8d��ֻ�(|�;Y �-�2Ŵ�� �县R�MpT�"��m8�[��s5C\2p$�2z<ɋk�|KO�7<�L�y��WC�c��ռ)��35�Y�v`��9ܟ3��,}z�,�2�9do�h8��ޔAB�WW�Z��̒D�&֏���6�tݘ�)h�^�L��`���_�rj��b�Qěu������8�'��&�Y�]WA��k���%a9�Z:�d|�lb�=l5�s\��i�o�����C�&nq٭#���R��������lA�O.f���E�y�ͤƥ��d�/wU���pG�SR�_�F1`Lxn�����2d�S�W��iU�z�]�cۇ5	ʥ��ŵ<��1��!>4�(������a�Uҹ����1���ԃ�i�urwI�>�A���*����D��K0����?J��L��aT�z����tT§C@~��%H�bu{-�<aۡ������������j��\����i`�e�2�h�1��MxY�߷�\p(A5��l��&���#��c��QcB���Y4핗S�
X5 ���f���]�%h�D�	n���d�N���B�G��5kWnz����3/]��
Ô,� �1��@'
/�6ȝ���l�nM�%�@��D���%	���%�Y"㚍�W;�[���q��ug�Y�~�5F)����TU���52��Č������1,=��~~R0-Ie/�b�oK���I�
����f�ѱJ�ў�ٷs��8#�b�\C�^ˋ���[��\��&������Xs�E�|��le\���Lv��ߏ�"��9a��,�+-4W�jߧ���ɲ��l�H,'����< �ԌR'?LU4Q������s'ZE��	"t���v��dy^7�f�=��wڃo�.���X���7��ag���z6eI��)��8���փ�]��[h������H'(n�Zt���ZF[`����������(��DO�����s�`2��M����ً �N��`���|�r{��x���Àë�2k�`2|�ϳU���������g�	�:ϲ#��!M��^S`V�=��![�GB#�:�����{���N�����0/��
���}���as�=B�|)�ur����hAC\R�UM�#�<�J���<�������},��k�
RI�����1����	��y.ޜ�@���~N�A�Qs�ԇ��ti
���Tų����}� ��-��G>�7�Z[����ՠ����������<�+<d'�%����SoZ�`_=�)�
]�,`�OC��l��L��VO|��u�� �u��`v%�K��)�� S3L߃���d���ɏ�� c�@���x��9�&/Kr�|���Eh�	�L"���+۫�K8\��0-��DH�!^�*mk���ڰ�n\��\����{mef����ŝ.�<��$�N����ay2�u�����f�Di@Y|zOI�E�%�����qDJƐ�Z{?�����Ѝ���o����c�X��vs[x	��>}B��9,'TH��3`��{�i^�F�⣚y������pG|n�K�X���T�b	�'4�f��\��U������# ��&~������o���dg/�E.�\�!������n�+��:ʟUѣ]�
�jp)�VJ����}��<O�ey�[� �C������R>�����I@�&�_�C�3���ϲ����=�����'⊱
�V�X�r{TO���O�/�<v��v��Q���8	�	����G�i$�Ij2����hc�Vem�^�{){�O��W��0ώ�������K߹H*ԝ���B�"1z
�MKEW���D�i��w�T��ڰ*B�,��]�7���1�&�u�hI�X�@���l�q[���R`V������eM�~�\	��Zhvt���v,���N=�#��&�D���o�EĔ+�fG���-'����j417\�̋�UWfK*c�+��q���LT����	�Z���eO&������M�o�L�q4�+�ֶ���5�����4�4�UO�.���b��i�+��UZ)�+)��c:�f�%*��U�vMd��Nb���ם��I�P�] ^�\��P<��K�#����.���ұdH�	xN���/Io��-�φX��#oU[���<���x��1ƞ]�8�B�x5U��"UQ��@ED��\�}n���L|���h�hU�zQ9f[+��x�'`�̂QIR�fN��ߴ�DF���ߚ�ڂT?A��hX�%;�#���ީ��"�� 8�MʅI�`qn���S1n�A@��r�sf:a���'�,J�0s��{ސ��Z5�W+����ku��A�[�eʟc�cVtAUN��!V��3Y��""��<��2I%ၖ}Ⱦ���4�p�"w�H��t>��!X�"~N7�O� K�3N�x�I��Ċ���f�|�B3zYöK;H�3��ff�^E^�#�_��d��{�I�S$c,
 ���!���m5�O�;�1a�w�ׁ wu�QP�*$�ɾE-<��&/j�u� �!�9n)�P5����=\DC�󟙘�3�;N_�^o�Ϸx��DP�G-S4����C �؆���S�X���#���Fu/��p���ڗ�K���ݗ2����)*?*�~�O���ƈ���؞�7K�y��錔�eV�?�>t�m�|��QiZۑ�樤*�<z��I��װD��k�YS��v5دȜ��d�l��ײ�׏�]�z��s�Np`�eӢ<��,�	�,�Kg}�O�I��3��:yd���]��y~}u�į�O���n1b���`�@�|�����"sl��R��^r|{�O������`\=%L���j����`$�W��O^��2��p>r�PU�G�3��.��^�w���́>	6w '�C��G�؀I��K�"�������Se�7u)q��R��p�W"�^�N'��-욯3zݲ���x�@%q[ɽ�z��2���e>ɉwo���.�̯0DL�'f2����BuҾ�wI�;杯����jv��UZ����Rԉ�Z�c"o��/�e��!��}z����6�;�Op�9V2%A�&��m�*-`�ۀ������T����)#������҆u��k!'�O��B�M�3qp�a�ǣ �J8׊��̠��0�&�iO&6�?��TJ<#�J�U�(� �G��S�cν�c�7�^�I1C�~��2��>�]����K�g�mݮl��C����RO2�8��S'��@�dL�EX�/5Z ���L� �qF~tϥ-m���;6��:�3��d4ҷA@-�=6�b�V(7��(�%J���Ѩ�%�+{���
�R���Wf�B�8��|gc�R�xGT����k�.J���[��6�T[��B�6��'-���)�0	�/�Q��0E#w�D�b�*��s��	~�)�o7F���I�wX$�<���cf`����]3t�}1��^�O�ÄGY��t_��ͯ�������ڸ�}= -��~�cd(۩Ɔ���L��p�V��uvJ4]�{�bz�����G�����[�H��u#r��R�CH>�?�8��4���I{�C�r�=W�5U'�KI_��J�UR�������V���j���[G-�Sq�be��j�Wd4?�#���*��B��IѾ��R�����ʆ>H�����l�$Io�0@���� �WfDe���a�!N�.ڎ|U�����6Hra��9�X�6�B�{{�,��Ŵ���Ȅ
e����bG ��i˝��3h�_?*�-�H � vɸ���5`�Q1�L����e������h+�s��D�9`�����3�\���^��)j-t���k����0��\I�,)�v��P�}��:�!p!��]��J�p�Y�-�Q��6���P�ѫ�Ϝ�t3�����V>Mj�{�(�L����>�ի��Hܛ��a���2�����	�2yF���	�������!��]��h+&�K��Y�-�����C����K�~��}���v��͐���A���������Ţ{<l��`�{j��$�v�
�}|AJo11\��3������?e�2��Ԭ�_��8H��5B�����Tے�ll� �a2�K�y������zZ��a8�,�-^˒E���ѹ��v�6��D&k����� ���o]V��z"���� R:������鶌����u����qf�<+�7c�t��N��>���PV������f�	��9����tL!
-�t�\N�BL��4_+��Y0���%��e(eDד�$gs���/2Yꋯ��,��	ph-r銩�d���� aoc۩D	�W�L_t	e����앆,��y]�_�����vus�D��YJ@�l_���e_�v��oF��Q9[��Z{��ψ�i���e`d����#�>H�le:����?����=΀���L�ٮ+ꤛ�1��S�����W}}����^-��z�S���Q�@%sE��o,����ڞŃ�b.��\�f��(r��pc��N/��~����`�q �<尰�h�Hw_�2������&SwDD�^;]cI���OH[�m����;�!?�H>3��Ԧc9���ύ�lM˜�Sj����;�w����M]Q�ޯ[��w�D��؅�ѭA$,>�ᘟT�6.3�EfH聘�;�����︿�7ɋ9�E|�"|k?6�A�L?�p��:��~�(����� &�~�����(���d��UO3�")�دX
6w"��V@��
r�GH���������]����&V�_x������$!�#��gŦ�!�<�KAP�A[:ؐ���0�	�GC�a���(��q��\�b��� ^v)��T���Gg��^Jh������3��!m_Y���D<��������!� ��'J
���T��L3[�i�/��O���>���^��\%�%��m-�{zC6��:����#���{"^�t��pN�^���-�c�����N�����K��[�i���>�����?G��Ǣ�"Wm�Éz�GR�,�je�S�c�U�K�u���p{tMpE@󣴦F{b�����}�tLC1C'�\e�i��Y{�ܸ���qP����չV�/y�Ơ���7^��+2b"q��&�E�r],J[nh�9)��i�v�����,�9H����r�;�&�71����Qy��4S��Pu[��'��ﲵ,�\����s�($L$u���6�,����8�ddb�Ǹ�i&"G�q%.xh
�_M(�\l��5Ϸ��X^����6�� ����&�م��1��7��~i''DUGP�ɺJ
]՘��]mpL(���]w�_n7B4n{'O����R> 㜹�48N=���.1��c� k�WH�ꤛ�����B7�%���8�֌)x�1��r���Ӗ�k:W�7ig����q�)�"�1��dz�v�{��^���^ITKz�@e�╄�	?Ķ\�P�&��`*�l-��*Â$P�E4+a�l:.��]��6�	�u�*��v�Y	�jp�u(c��g��@��^\���֬��Õ���{��Z/`ߕ��_��G޲��t[����c���{���y#�%�f�虋�_��V/��2V��V�K%Da��W�^�PRő�ނ��lI��-���S�;U�P��3�Cm���>Z�W"��t�<�j��CЎ�wr�`����H�{��>��m�t�{V�0&�)�F|�����Ҿ�`S�o!l�pD�*�SǗuyg`�ɑc�r��<�yd0	��wd����96���?헥�#��r
�k�l����@d1���%89��]-#���!Տ��OR�ƎCRpL̸a���|E�#��&�~� ~�s�C�n�!:�K�~�FKHu>��E�s���ςKoeP��Og��a <�G�� �1�H��t����z�%����P��65��&�5����(�ǭ=�zg8���l/����OE�se5e���I��j�#ǙL�[ga��\���#k_�x-�I7Y�*�XFi�A�d�=�-��B�bb7Q�>�4;����8�D�\��FENq�t��F��_�
]�c����]��1�r��6�b����o�>�V*�E7��cU����d�E��a�.,:��A�`��tN*ɣ^m���iz�e�\L����i�o����g�� �� ������$�'¨����؅_Z9~�;�l]u�$#4�Բ!?���N��:�;�>��KL���g֞h����ߴ��N�%C���=p!�^F�3�h\�ݠb�h�t�~/�^��������L$�����F@O��0�����*��͈��9��be��  K��ީ���th�t�#�C������b6f���5�:�Fy��ĕ���-:�� �y��偧qg/t���B���	Uݥ�4�Z!U��w�=Iػ����pJ�U7@�����^��"y��k�C�ܵU��B�@k3�׷>���El��b�����-���_g�3T�N�N��*�i���|O�Cѵ�$���\]ta>^<��G�T�!
�#��U�3�R�ر%$�����>�E~�����f7i���.��%���Q��h����!���@q�F�G�S�<�v�c�"~ku���VK�2�g�Ǩ6�κ�L>��g��7i���2H,��������û�`�&H�Y/m5D�q�,2:��ʩEr^(�q^��H̄�s�[,e� ,���ߺ�4���� ��/Y*���/�,���gEŪ�~Q����⫱$K�ҁ��=�������t�b��F�+֩T�sJ'M���I�a�9eǀ8�x7L�#wygA�zg�hԴ*BjXൄ݈�DM�Մ��AeEx�����?��K�>��3w5������9����T�[�'̻�G9i�o����)D<!�]�ׅ,Ole9��G��~#7��v��ǖϕ�m36����i���;��y�]���vnO:�����������&F�,'�8U����d��d��z��f�n�~�Y��O�u�#"�|q�b��0ŰK؈�ҷ,y�Iy+D�!��l9�֓Sڸp�t+��c���\Ӝ��^J4���	=AW���U5�?��L4ƅ]�����UA�kV�$o��ۧ��K��fT���y+"|0��J�`�!~�c��OɃ�4s���4v(�P&�τ.�z�ٓ�Z�y�F[�,�J�G�����f�f�".�]��4�p��w��[���茓���])*�����G��	�]� )��`��m�I�/�TiMe��N��c����!}���=�W���Bh��(�A���m狍5S�)�"�A"���$i�4�8�6����(��m��{�m����I9���(c��<���@��:G�GzI쬪�� o-���#���|��U���Uo�Ur��S�+�(�	M2n���Y��qx�����G�	�]�W���衮_VMZ7zz�Oj�;&�T9�`8g8t'��K�Qˁ�"#&p�	/�"��<bA��{ �m���Y�v+�SGϿn��/y"�_�>�d�I�9 �f���r��c%��K8Y���X�!�����:("��i-���ܿ�S=��{�oF:����6k������NK���Y�Pӧ��Q3?;��p[�B�6e�Z��m��0�"s�tt�X�䄧���N��y.`�x��?\�����(��^�X���X����(i�9���E�˪�4�_Oi>�m�0�����{��Q��`#y~�;���{���.��Q��Ш�d�%Ŋ����_�����"'N�����V��-Qg�+;C�̦'�b�dG;���^�WozJ;�O!k�?�$a�e�I`�&e���4Z��Ty�ѻ�7palQ�*��P롱.ǒT̕��I�4,�9�CF�U�����@�#IǼ����4©aԂ�r{XΓH����p/v��cWQ�h�"����`�~M؂k��\��%����Z��y���Z��R�ON6�Vk�q}�W�B�M5�lg���>�g�n�󦶴/�/o��)���������WpI�臷ks{~��{�S�9m�R�=����� �E����g�=�C�y�pfŎ��'�fb�gR+-���z��_ZǓY<��:N�E��!��Z]<�x��^��jfI7=��0�#D���m��iv)�g�L�d87�c��x������q�V>Y�a۬ ��(`�]��0�6���xJp'����o�[^K����3��}�j%�uݫo:N���y&�\X�Qt&��rK�/r@#�)P/D�Fopgw!j((�Q=��Q�Q��YZ�j�Ӡ���C�(���� �q:��ԝ�O�A�ulkD��[�,�H���YA.����HpG�z�x��:.��"J ��ɜi�����o��_�9<�]�AՋ�{�M���Ĩ���b^�Mq��|��S����2�Hf*@��=7�K��Y�Tʿ(��͍ETӾ�=�&UO
 �4����{ޙGX�
5����f��Y�����F�D���u?����j���n��������w���)1[E��ib}����j�Rk��6�f�c^QH��%u���%m/��.�z�g�Èr�N<I=ɬ���"w���I����n�m���x�X��c3��Q�J������-ds���g���4l���B�59�*(-�����1����!j������}�;[���u�
~�Ɣ�fcᆁ#���6p�J����)����b���H'�_�Ϯ�"�04|�T#%q�M���.�Gz�ur��e!�,�1�G�hF,�c�B9�#P�ld-V91*�� ք���."�I��!鹈�ېv�{����K�=���"]��I"�J ޿G�	�'�aO�JVV�FA���f�M+�	s��P�))�9y�ɖ�f���m
8�_��:e���*�s>��#��/=|�|����:�
��w�mn���r�����Q��`��f�Y����f�~�n�&�S����ъ�Ib� ^�gI��F�hj��bk���Cq��d�Vɸui�=�I���?K:��y@~3��x�f��Y�'���|;	�F��g�k���dr=�����xZX�V�����d��k<�V��P�s"�Ɛ2Ԏ<H� ,���c������ZJ�Ѐd<���ߏ���Fo��gw{ft��y�Uh!�a;a0�cH��A���^]��x��,!R�WS�-�P��X���(��k]�"	�@w���ѧ;�"�2�����v�*�����@��N9U�m�W�5pl��\ֻ6�ȗ'�Q*;?�9R������9��y�2;Y@iW���ge�����:�8�cڨ �y	��p\}m�b��; �?���pO�}6D�~.&��H�j���+3Ñ3�N�Y�V��T���ߡ��>���D���!����:uF��腆�(�d�N�x�����̽�&��t쨉-�`n$:FDK��jK����6����=��c��l��0�-=��+�Y������>�`ģy��/�p�B�o�����d�}�-�z�?7�����M�n�́W=����������yꔐ\h��4_���B�T1��03����]|L�+�=���'b�"���L3�l��>ĳE��۲���]0S����q\fI��3˿�V�i4���o3�F]|ڰF8���eyoKt�����ƌ�&x
��"5pˀ��r��(������1{������.����H�Q��p�=�r._��R��D/�pW��ω�E<�c|������@|A-uG]��������kH�K4���T��3���wJf�lS���yh8RCܻ>Pu�a�v�)�_���Ǔ~�k��kx�6��?4�Q��!�#�j�Ոl�N�5�W�R�牝��Y6C^7�S�3��&�r5aZs>)���p� ���v�#(�ӊR�q��pj/@���e�`��*Sq��������l��]22ʋ����W9VQ�#W<Z������9P�w����Lɜ�����5�~�m�GV���z�pC`[b�NϏ��6H���x��E�[|)"��a�BA�?ό%@*�D�k�3-���웁���ȶp{�[6x�#����.m������ @j�e�TAc����4�e힘����0w�O�ى>1c���s��'_B�Qm�\{���+b���yK���<���8}5Tte�ʅ�vQ{��v	���:��	"�#�Wz��:��)�X-߼�1 �,�]D�ͨV(;O[�;崺�7��Ȥ�C��`�?ptb�N���������k[���K9_5�̂��f�� ���SmV�^Ě�w`�4��>e�_i��u���Uy���V?��ef�T�|Ϝvmp�Y���'�����CB����gbఁ �i֭zy�������h��\���e�� �B�i��]� ���B.���6��Vo��
T���S�\D���o/�k]W�#Cs��R-(�p-�2����Ώ�Pԥ��<u������*��L�J2��D�~�*�c7 �cY�8����1�D���L&���Ul��WaC� D���`���]t� ���Sm�,��q��|��O��/}��c�fO��nPSѐo�;(�N.$�e��ъ?�_�]�o�!���E&�d�;�ஜQT�XP�Bdr�W�s|H�� ;a_̑������N�����U��7~ܡ���5�&O�T_�_P5kG���m,����Ԯ|��v�ǅ�X�?'Y>����]#&�H�H�28�[�(��I��f���A�ڕ2��0Y�va!�kιc���Ea�J,'��|F�n�(߳�?(�D�x�B��3�b\�>P���sa��j̮^<�$�nl��� }f����YtAv#6�T���Y���JpT{��o�o���]��fok�]�CD�m��B��^�����ErPŅ�Ī;n8N@J`��ě70��!#�y�q� �V��S*�i�����\yG��綬���.�?�g"9gr�cq�����a��PTJ1b[�
>>=B�
���kH��l�R���$7���/�:��_JLȂ�+ߏ-�_a|F�z�GO��t�W��.uU��&�(����B��䡁
4�[��q`@��»�]�w�j�Ӿ�N�������{�$�HdoM�����p�[�l�����x!~���u�A s�	T�E@����!%�6���L�,�f�4�|g�QH�; � �"��d�B�(�%}2�m����(:����/��)j�UOpqR�^�@bkK}*Y:��X�x�h��2�]����+�<�iְ�7�p4��A�*E��Aӵ�������e@Nvg_9:���;����������[�	?p̆��<ٜ,��%�wm,����Q�B�'�F=��T��{oi+����v)֜�rZ����kE�:�H�S"��z�������:�S��,�����n'q���qT���j�d������Uvm�5 �)G1���5��О�Hf,����
��V�X�z��ܐ�@.�2��3�<^���q����xr�����Wn<�H+���ic���!�z���W�C�7:��1:�c�'_j_�>��b�z���K���,������T��d.�2�V�\=_���� �9��x0r^�(�LJI�����+�W4M�7�@������jYvyp���j�2�?7��]��:!�oeP[:f��2Mj[�M!E��m�~�]�0N�5��g��g(��Q��|��4�Ҋ,R���:~;։���т�Ye0c�BI�������I��5#e��X�L�l>�����@��;��a�o���hڢ����czx�ƪ?Yy�o�U	�|���f��7��<y�Y����?W.s� ���R�d����v{߀�k�zk�,+���wCb�J�����4t0��@`��!��6�?��؞iU�d>�s�;}[�$Q>e���H����#�΃��a�oz��V�.����6�{�aZavև $ٰ{o/���1��U�;:4٥V/r:7��kI�~�>*Ё���4��������n�oӷ��Ah �!q�to�y����Jc��Z>�[>L����di^BI��cS�$qq�o���w�:�'X��@��ɣ�5������Ch���ΈAe-������s���q�U�f�JJH�+����Nx�$���m�͆G<N03��O!Á��#̺��~����C�����]�?�M�L�~�C-�g�D�a�ft>W샫���k$QGv_�ˇY��L�]	�0�(�]���Ы��J>;��O�2^�o��\T�ɽ�^�)���e��?��3P��O�B�į���>��<��A]I���r��]��Z���3{C106����5l����f*s�#P�L��.�A]y�)�{l�$��٪�w�$��Z�{i�`��S��O�.�ݕ�7�-&�·�"��jV�v.P�s�j`��/�Z�ڃ��?Q���v��,�(N3>�\��N��0�sJ��}�� �����p���o�Ϻu�� n��B�M�\����/&�><�y,U�=�cĽ�f���<U
$�9ń�l��m]����3�P�l}&�k�q�KH�A�R�z������w�2:m��c�����S<�ɱ��-d`�����J���F}Qr�(>�W}��o��"k���6�	%��~��� �h��@�?�pC#O����C��jX\�-K�� �$��Z��zFRjZ�%nKF��x��_&�8���E�e�!4�a!�X�k�y.���ZU��ypW�5���:Yn�r��t|w�$_<Om�ϑ5� �'h�� �ڊ-�=	Sp)�#�˭7V-�$�n�q[�A���9`��zF�0�k�X���߈�G�����b��O�&.&y_�q�@�*�L���ͬ�O47����<���
�����A��V�%�	ʏ�H�s�(�p�\��6������Sk�^8�V����ESM�f~	F�j�������\�)�����`��ְo��n���k��e�E��/0�8� w���7��9�R|?=�D���_:��������r?�J�i����ڒB��S�r��v��� w�E�0z��Ųã��X}R:��NAΆ��L梽ZXՌ�0�GӉm�1Ջ����Ӫ"߀,[3]F�����vo:Ტ:�.� �͚}� vEt_SZR@ʩ&@%��2P��Q��z�D�B�u;��W+��|�`)k�1��A��
 a)
b�����[���e�uh. ��T�H�2�o��	���<�Z2S�o���c5
?.��C4N |Pþ��7�	�@�!f~�f4�dc��s=��r���g[��r�� <�V��/��w7���G�r^�����i�d�C����D��sbT2M�~%q6q�D7z18J���n�aL���e	D�H��L�g��X�1u�Zh#Y$�$�*)����Vd�u�Sˁ���$�x��:��Qc�~O�bF��%��B�0`��%�c��Y�A0��B*�.T?��+�C�o,�~{�;+*3dY,�>���;��kZ�A�a&-�B��M��"�Q��C&��+��Q��f�
�;l'xB���k�����]Zz@Y��^�Q�_�3�"��I��m��6^�T)�s~^�۬��;����"(8�T�n��]�[����� �ա��A4�#A�?ۈ�9r��T�!��<].��i�az�1���ЃB����_Wo��~K�:m��Uq����H7(O�t�&D�L��J@귴���X�YŭH���#��W�����N��6,�#<��0��1�I�f�Q��xs. �V݉�`p◚��4�n1%� U����!�_��F[
��E�8~�ʬ�T#�Y�B��or`j.�#ߑ�Eѳth92U�rn���
Z�����
'�.���D@��m�MF&��?����7��@�Hg�&7�|�1o�����VoP')L����h3����bĺ��T��nkKʞ!k`;8N���D%V��į�>ѧ��������f����&�:�Q2$������75��M�a�9n+`��;���ē�a��DtY(�#5���=5�QA,�雂[��v�k��o����x���bm�sN�����[�Q�9�~��7��C~CJNx<��b�3�Cg��oQ*��V�,D(���+Q�p� � ��DC���&1�UB�w�x"�� �Y�V�<1Z���F0)8Uj��X?Wk5l�r�6�k��ѧ��5���L����G��g9���IҺ����׏1�RHQѽ�n�������'�Juj�s}�hr ��L1��R�x�Ri&����Dϑ�K'W��������߳N&�ᇅ��'A������%O���i晇�d8�r`
d�5@��ÑGɲ�3r{��:xDi�	�lz4���Y{�O����C��^_��t5K߆��/28��0�<2�';�&���=G�'���[��/䁢
��G;g�z�� lT+A���wQ
��D�Ӌ���-Mg�H�\�Q@�L���!a�R-����+�7�d��W�_����Bx���9Ԓ���7������Ҕ3����4���ŷ�j��2L1,�m;l�ewDj�搋�r�|�,|��d��?��{���Q%��S���B��4�w��/�ZSm|��Vo}��pz�v �\�jt!�d-�n^=�1�)�����ru�|��/%���U�Y7�ͦ�{08���0Ѵ�#�ߝg���Wf�a���ۛ���ʐ�����.�*�nH������հ���l�N~���l�O����.��if\*���K�LfEd�yHo����Q�q�y���b��� ��$��s2�xxH6fך�'���@�2�)��߈'����a6{��z��6.V)jh�{���� 훔=W	A�{��͓��m�������!e��H�>�ͳ�H�c�R~(���<�ռA�_g-'�<4��e�lǕ�`�]8I��^��i?�o�&/i����B���ND#�NT����AE�d�C���O���v���ؒ�ԯ��(�H'����'���,��dGGd��o���?�,m���h�n�����fD�-o����e�M�>�c�)�_( �AI���z�^�7��������7���2dC�~��1q�gG/��O ���-W���K���o�5;��c8z�(����=|筊Jd�Zҹ 5��@�M���x%{P���鏱�w?��A��M��G�ޥ)���)�B������U�q�����3��n��M`QM�ʠ��jB�g�bʇ^w���7_���g�lĶs��2��sc�
�C�g��6����b]��aH1s�8\����	�ܷ��k�B�Ƽ<3�Ȏ��hJ���&},��*pKAEⱢ�_���S�я���y�(�@�;:<��5�k�V�۔ƫn:�P�8�����͡pa�p��poɹ�4B
�c���|�X�_j��e]#�v�
5E�<v�{F3��T�l�I(�Z[��#�!��@##u;J9.�A�}�*�z^Ҏ���ℚ��dtG+����J#)��oyZ�by�����E� ��Fs��ЯE�Whe2����h�2������ہ^7�J"�����5%����6�1As��&�45�u!�ľb,#�2T��{�B$l9�����k�f���`@��wQ=�����NíV�/�yӪ8��z@,D��l��AJ�{O#�l�;.]�D��f���oc�%l��BFW���7�A���
�臯ؽ$���\���԰�E�� U�\�Л��~}��ݩ9=��M��%)�	�/��_�������l�������Vs�ă�97Th��Ʌ���R�9Y$>6k�0��d{)��a�˕v�o�V�z����a�Y��9�ٌ����ܼ��<�pLG�J&�,�
e��(@�Ȥ%��-(���WPj�p�Ç�Ƥ�n������)OXϳh�RK6
%s��f�~5��b�9���2֝-��v��ռ;�uݿ^��rC���
��� �����E�.��x8��Oh?>��vJn�g �l-6+.,���pt����0��ۤ��y�Xk��U����<�%��N�<&���X�_u�q��7r|������EG0�Ga�b0�s ��2�"j��9�9V�����E�,�@ץ��=�|o#��xR��#�-���U7��Ҕ��*�l*�Qk'؃I����liM�]*�(<�J
�̍~�#6$���)����ޚq�)NW�"֔ә�ӏ~4�_�G;r�;%b�I?�G�ْ_g�ח{wo/į�q=������V�VG>�|k�9,�%J��$��K�ȧ�;p���ß���%�?�Bx�����\Z@��࿺[Y�i���W�6�9�P;�d�c���=
��@p�<F����>^�U��WT��G��[H�yF���8�d�H�i^�݆�:y�"�"���r �X�Y֪���j�	��A���ADT�4����#�-���\��Ҏ�o=щZ��(j� �<$E?6iрU��U�ll簹�뒭�FV�b��i��� ��#/J�y!_�56�!��Ϧ��[Nx��2~��0HV�˛�)F�Wi�7�����lJ._��5{�#�<�73v�9�B"gъ�|ȷ��^��&Gj���t��� /{G���d��h�Z�@�,�n�������ӢP�ʪ�K��.�=�k�FyOv�?����t�i�HFM|Kr"H��e��44�oo�E.x�?jn&(�B@��󵛃	����/�IevKL�`jU��
L�Ճ�6\��9��R'/^������(���B<�}�����-q8i�UMexp��z:C�$TZ�j��a����W�'n!�����Ni{1�ZA�k��y�8wvC��P����d(E�V���%�rQ�������t��������l5��-�A�(�fG�}0�f��⻤���ր��@
����C"fUj���K',U�	���B��n��W+��~Y��UB�mi1��/I;��Q�ޕ*0R�p���:�o�";��k�$�2���:.�Is(�ǚ�p	�#�� �b����v�_D��D�}\�L��Y�4�&���6{�s��ݠQFON��g)��hTl´S���lV~�M,js���KW\5ۊ��;d\̺�)�����0���G�;���e��?�2����"4q��Sqab��l�3��o��C�5�s�&?���ì�*x�F(�3�2�i���E&���0K]\˛�$6޻�#Qs�LM��ؿ�n��x�w��3�%��?�j��ѷ<�H��5���[�G��H�/]�QC�^M���.�����?Ƣn����m������Ҁ`�����{%e.�����ea+8���fw��j�=)�5z
�_|opƜy�5�?p:L�oa1���*W��8�1ն%��}�űʲ��UYтZ�<�[���J\3��
J+0�����+��<Y����~k0�3qG�zUt=�<���3����^�-��:٠��f�%���xL!���4�	� %����gSVkC�$�q!bw	,N��G���P�X &�q��|�
 v�Ց�y�'	��3������\�?�k��#@�Y/�Z���Ҵ����z7�$(�l��>���#�w�~��w�E�����\�n,�4����y�%V�*$��{��;h�Z��˰p�U'��"s��$tK��՛eU�����؅O��!��x �ۨ��_{��d�ou����Cbc���ӱC��c$'��hZ��tC��Yh��7�fp��Q�E�N��p����R������Dq��^<���{�Ə��C.
pc��Kõ�p��|;F��o:�	�����!k��s�ɯ�ÃN2TĻja�n��ׄ���l�ނ9�`�s���`��a�N��G�[�6�`��.I�Y��~M�8�$����6����KsC�������Z�%�s��JW������+7�'��ܕ%�*Jf�`m8D��r��4�2��y�I�L#ó���IjlP��8굩0�Ϛ�,3<��%�/*�6�V��O�ôzz]��c7OA���5��>,>O56� ��X���#���\eYw��K`*&��D4�I�y��%̎S����+/�;��upu�f gD�y�-]�rX����*���jʃ�8�S�R���,q���	�+��#�n�6.huj�sJ� f��뢟/#U^�P�3-*�q�v�0#��(��׫~7b.
gtU�	���R7'0<��/Ӳ���62�KbV��7��ψ�q�����@����$���E�9���=�_�J��Ϟ��Q�e�#J�:"�G@'��F� d]z!�(u y���V�,hF�JT���2��mK���ZQ���G����y�0�ȣ�i�H�K�t�n2\FC���P:F�X�!D�Z��?�w�d�-X��jw��q%=M�mڈ�N�h��VmZ�Ҿ�x�p��v������ϰn��
$��B�6��$�$��g�a�d3��P���T��W�{~��42wC�5;�d��Z�/����) ���˦)�奧��je|�~Gn��VI>Ѵsg�<� ����9�s4�Nx)=tX(������	���8�f1��F�1�H��9��8����M�%�;�F�!MT<��,(NZ��X�z�(Y����ĔK�37��U��[��\p.��.p�ԗ���P5Y�M�F/�z�30�j�1�bl��һ�,RrV�8�]ѐ:G�$T��ntP�Ԥ�ekߪ�=��ɀ�m��V���B0}c�_���IL�E��⃷��U�����RO^��AG�o��v���g� 2X;��mȑܜ��/`�@�s$+[m�ꇋT+�u��kj�x�O�xwR��(��h�D0��(�����k�#�"��9@�j��=�,~���6)1O��� �d���8�;;Y���y� zU�������ygʵ�C���r��ҡb=6�יW�K��/��o��x7�-wN��Hч��W�ki��3{*lʿ��}jL����1R�	��ۇ���! ���1,˳�pN�E�E����Cn�G_�4q:�������5T"3&e�櫟h�c*�2��� ��2�$�{����ڇϟ�.���#ث?#��`���%����~����|�,r)�S�}W]�>�$~MID��j̭��}
.��:���U�-O�8�/�~*;�(�wHI��B��޸! �o4���ra	�
���t�҇�aΈ8:��u@�2Q�_��F�D�:JW��(��{�U[�H��
�ZŃ�)^�v-�؈9�Lf4�:��*T+�F�jA.�4����VczZ)#�׽Z}�Y�;3���t��N��6��f7\�P=?������r�4DK��U��5��THZR��]���8k��	͉�����w���4�;��$��:�Q��LS2{
 ��йx����OL2��i(�^��EU:���r�H��VO��(\r����lG��s·��%�d&wXU���V��ă�ղq�W}����ڷf�� -��.UmX�H�? �G���h�?��|��*�"Y��H��Hz�/��}�w�?��A���`�K A?�� ���`�(XV:�l/�ZF�~wͷ�c	S�ބ��uN{���Wj���k��O�@^��w^��j�7�XD�ZÀ�>��!W�7*�)�w�(ϊ �a�Ԙ��ϑ��E��Nj9���,�Kh�!O����1$�Xe�˸<�S�$b��?!���Paح���bMR���(��D_���sͣ� ΖG!Tc)�ݺ�+r�v�^��u\v�(�j��r{P�Y7��U���c�ΐ~8�Ј} �m��*��b�嵐�&�U݉��u��]=��$~]j��A�����o�M�.��7c!XĆ㿡q��}�s��[�e�hdM���Q�	�K�R�5�ݣI1�Wm�M�C��9�ze�5�.C\����d��|��\GL\x���Zt�W��!l\�]�hh~�\L��%��M뙑jU�X˓<X��{��7H���&�:f7���'3:]�S��LM��FRϢ2V ����
}$�\Ӥr�� o���](� _gD%rg�KU��D�ߒ�L�.9|�hFaO��~�&ۣp��x��O�,O��NP�R��[m�� nr�(��(ZՑ�u����=q�{�Ռ��:En�MuūXYK�$�]���\� ��H�7ƭ�>ý �[����"?;-�.�5�Լa��n�<�<X_�����e'=XRW\xf$!a=�y�,�l��DE���a��������C�!ч2J�U:N����2�+��շCA���O<� sA�!�lp�E�tp{�%��N�؃ܑ/@���x~���$����G�.ŧ:V�7�!�m,����E;���?<>�e����b%f)5�ё́�����QV�ƙ�`�K{�1ǈ������ ��y�f~�b����e!# �7#���\p��R!ϏƊ�|�xz�ʾywNaÊ����=.&�!V��#o@��I(`�T�7
���8��~ZFb��5 '�)�+_�E�H�:���h!G�$w]�����R�z�C�M鯻���cN{�z$HQC�0Y1	�_�M�_Qhԯ��`�+ͺ?���݄|�:�K}UL�\��*�z�&��]8o>}0$�P��T� K�����'ZK*�1��%5p���T�}�;W��j�8g��O�Ux �L�:���o��o�
ē��J9�UEY��s�ܷ��q��b%X�뽁%\������j>zY�5���V�n�λ�<Ž*�w�7r��G+]�jbY���^�UO|K�8����(����F���EB3�m��-�}'ys��% i[�j��+�4��5F��Mf�M�Z�(��i�ܙ4Iս�F�KGbģ=Io|ɯ �3��Z{@a����W���­�1˧��5T䞤���-Kv���ʌ����"���*��,����]�~�B�̨a�O�9G�O1��X��D���u�?�A�)3w������D��п���G\N����Ub6���,�;��z3Ã�	n	XBH����ܔ����o�ȃ�$�*r��:Cv��KG�%�o�hٓ!����j���H�01�g�	�<�Q�WI�ԒC�V�>�SX`I��	T4厂�p�H��v�&��S*`�(�г[Sȃ�4z���N�$&)$�޳M�=��Uc�%K]螇��%�Ԍgǣ�T�r
�"��4.���m]&Rgc��R ��[EN�H�
�D��kID�9�}y���d��H�m�����������&�+e�dY�ӛ����@*�XKnA �2��6��.%�'�L!l�3g��j�V�J���d�����JXon��=�m��<�D.�^Sq���c�!�灁����Dd*EZjf��5Z�M�חy'�R�&����l�J���ɗ����lp��b�����V9v�DP�9��=�\�ڿ<���A�a�g�k����?�vHp0�sɰ˼�g ��*�t{���V>�����.�kq#�n������"�'��\��#)���pD���Na_嬈�c��{���x�Y�*�xK�����`��Le�h޹�P�Z+��@ܲsk��+��q����$88��2x�����NS�oe�yuFI�{�-e���+W�ߗ�֖M�����G7S���oR���bʙ��k�<-9�
S��f�9���v�3����HhrHژ��Jw�y?�_,�VN��-Y�w�M�czײC�>�[e�L�q��Q�!_�4l	q�(_�-�m
�wS]�(��}��@�c8��o�,�a���a��~���*���K, |�n�AJFN�X�|�F|� M��V�_j�8�w3]M�ߚK�iyR�;SY�Й�Bja�M�RZ��^{cX3���^�_s�����"]2��P⿶��7I��8�èoP1���q��a��5)Щd-k��"ӽ�7�6<,��[���C�ޟ�xc��Lc�cg��k�i��xo�y;��[��-k�>��[A�z|/�4*��j���-A)VR���7O�I��O:�ex}�^�����Я�y�$���x��]��U�"
��K���(���1�Zvj�%|�_^�JZ-�!n��B�����W��J->�(�[^V�/}N��|Ƞ\Un��`8@.$��褘Y�j(�^���:�%Sf�����6Y��W��8�L�RI*��υ���+ʃ�0�9��y�Ż�@�~(�m�צsaķ���:���o��3��}QqQB����1sU�������ס�2ОF����ʪ&�	�����e�yˀҠ�
�-Μ�����B��:K�m,���l�}!�)�vj!��T�C6�wQIyK�%b6�U;!&Z�Ii�����[Q`[�9t��Ak�O)�XD���F�N�8�;W6�=�mB�.�s)�$�5�a�j�'���׋��3R�<�'Y�;wk���^(9m�wHX�f�Y�e�F��X��(&��Ynf�����\.���F����w�xEn3-�e��}��Լ�ĉ~ ��"�ߋ��ps���c2}�����]f2L����8�D�j�ĩ]*~�T���L(�#�& ��5M]5p=������fC�e���h ˆX����z��д����e��P��o���؁�48ϊJ��Y������e��pP�)�I�B�������3Ga3��zh�c.�%<?�Ӂ@ufb�	�+)���҉H0�,t�ᛈ�$��L՟b2�&��� ��lt�Kտ0�y�F�1��!�Xթ���aj�oU�t�A���I�a���w4o�9=��t.����0�|Wh�ʩ�I��Hf�>!�{�(�������8�A:O:P����-��x��8Yn�~8�F��������+DU����K�������Um��
S�(+��AS���ء�6,&�! ����ݵ=�9qO���W�ཨ��B*(W��'�faN�U��4zqz�"z�k��B�UM҄��w�B"�ѐ.�*D-�d3F��ε�����PÚ�Q�0��v]�#0zdeq��d����38�R�J8c�bZ��}�8s�2IًL��~�R}�djk�.���]@�G�+�X<I3`O�0P�yɃ&]
L`7�#<5���q!c�<aEz���T9	Q�$&�T��	�d�&��[��:$� �oM�[�]a����g稫r�;.S�n@�p�?��Dnx�_R�8G%��!�`�{�PFp!u���h
1)G����)_+�
[�Z��Įn�.]={�Z�m�	�����0ߐ�X�q��A8Vp���|�(�ī��R��p ]$��_~J"�T�����SzD�����>n�|���q7�H��x�&f���/Y�?��V)y~��}�;`Ԩ1�3�7�n�ڬX�u�Q������Lx0���;/�Uk���[F�s���xP~w{ͧچ �;]Z[K9�pt��B':���$�z��� �:P&���"I.�h#�����fn��Y���-"�i�@a�,}-��9n���}�L�v�b�p�X�V�&AB�#x���	;	�r�� ߴr8�[@_����"&�Z�� }p4� ��6�D�������L1�?���Q��ۘ�c�n��ш.����9V��Tx�ҿEGv��m��l1{[j��Eq�!]�^��Ki���/B��5��&�|e�Ŕ���M��n&��/�}���|��ƍm�Q�/pv�������O���i9Z�kX���e��rl�w�X���KH��l^�U����)?۳棱�&�l=���.P�f�g��K�����bI����� LUV�y�S��L�^g7+�U�u'q��TT��w���7m-�PJ��&(�{�<�iu�+��Zn�&�����6, ��$=6 [����vJ(g�\�eۤ
��+9^�/�):Ռ�~�6F�j�y 6�B���K���>E�P�N Ia
�'?�`7����:"?�&&�W�wZ�V*�;%s�D�Ϸ���7Y�l%�*�E�wѻ�fY<���m��ss�����	��v�i���`"�u�A�)=(E�\[tS�����Sہ�x>$ �VwU��1��CZ"#�����N����-��2��a������6�G�a�N_�8�׵w<��ͼ����^N���g�L���� �>N�ȲE�Y�<R���E���F�J�����lۚ�����E�8���An%ZΛ"�3g��ʶ�K��Z�6��HOW��b�����Yn �}:�vly!��(��:K68����Z2Xv�e��������)L�Z�.�k�z�6yKo���Hx�Ew�y�#m���D������3!��4��[�֬�{B�r�<յ@���������n������}��Õ�`twy��qyF���|��\(�L�f��(�?
��ߕ��r��ч>]��T8���G�AOV������2� HQ�g���7�	~v2�f�?M��w�؝o&&MܹH�
({����0)�V��DR`1�""g��0^��v
u�.�����tV۵6QQ�#������12�W�]�g������F���#S���tiM�:���A�m�ￇ�޴�R�j�!�����*垭I-�� ��A�q9�.W�@���	C���j!�2WQr!^~�*̇wd3̐Ǽ/�����_��h�W
���<;F����o�H"@"����.i� ��M9�1�5�x��>e�T���B����vE�W��<�0�Qs�����F��4�L��@v߲�"5�3@4V��0��1�i�~�r�@UoO��������r>�S�X���dLx��Z|	�7�#
�t�䍞l�<�S����8�,��Y�+���v��L���Kť��L�6�����rb�)�xm`L͘�N2v�F�UO�+�Gfլ� Pm(�rD�b�GȺH���@���F���Wx����j ���^6�m��c�n�"-��<V�rZ˰�}��(�uDT��۞�׵�76��UlY�>�j�<�̐�/�!$�&՚g|$�O�}f��M߸M%������/bp���^�t�fVS���?V��W���c]sP90=�~'k�q8�j���.d޹�G޾���'3�L0!+�A��.,��1��MPB�~� �� �b�#���̀xy7�/iEؿ���n��M�r!f������
�+�b��@X���T�!��|y��F�0 �ss��07�?�E9�"}��8U�g�)�H8�t$#�7�"}B���ܘ�}��,�s���zZ;`����r?�*�a��)?&ځ�����n2��;��Oz��6/�2��6 A�W����F�.�a�uX�����p���Ψ�D]��z"��ъ����S)��1\ǆO��c
NV�~<���b[	�����ux4��^�(f~V�S��dS���u]�ߴ��h�۬(� ��6�ȓ��ΰ�};�F��I)�����hh��@H��GH����۲�?^�����z�F%v�cGݎOM4.�� �N��d���U���Ob�CX ��m��.A䠀� ���֐��׳c���i�dM�E�~��0�$�fT }�47[L��8�- @�U a���7�L�����Z3'&y~�#ryRH2�|�����*�?�cP�Q�j�$5}4�x�	kś��h �S{�qќ&�W��=6~�O�F������@������h7(���c�(O-��w��.N�Q
�WRjq�.΂�Z�ߞ��8v�5$�]�V�����]<�~��:H,�k$���dLԐ�hF���p��q�K��b�� �����nv=�1�O\��>)�x�5�2�/bށ+2ߘ���JL�����_~t+��������D����.X�2������1X�u�l\���艊�|��R�T͒�����M�s�G0��YK�;Q�����`� �~��0�Y#��Eb$#������W
���TE�q�f��ٛ��日�2LtL)R`fr��?v4!r1�mf����p	ɓ
�C�Xz�T
q�8�h���!�� '���H�V����4,�:f��5�tA_�- �O+���(y�,���̟/�v����I�C_Ga���x+Ǐ�"�����B#�E�3�K�JB+���!�zܠ�yd�C�'�F��a3�RIkT� �G[�/>x�$X\�S?\��ѥ�h�^*J�ߊ�"�{ҏ@��4�M��@3ӯ�i��;��-���`�* ��a���D�_��?Lo(MwZ�1^�+)7�����'c�]j���y<�~g�MF��L�:/��U$�-7�La��Z_B$�t-]�ˢ��� 8/�@��%MZ�X�w��O����<dV{ �2�X��	�������t����R9p�&�^l�C��Y�n��4&(G�;�+>����ޜzFt4#���������5��OÄ�e�.����=�j��2�ھ�3��+�Z����	.��5Hj�㝽I�p%���W.��kX�~%u.G#����:g�M���at�vZ�nշ�����m��[�-��V��Q��T��|�
@����F����p�BṄ��TD��g��*K�"� ��L�~#�l�րp������U�1���P����T�2,���5�,��r���r�FoD��U�̘Tw���4�-�~�p�� E�ǀ���?��z�1H�l�J�Zǎ��f~:���̟ ��^��ؠZ�q�H���-�E���1o���k+L�~�p����>�|E-[�!8 )����@?$�9�@�JI�#*���z�5�M3��.��Z�O�Ψ	�0W���7`��eȸ��_b�ē�b��sԕ!��C������S�X�;,��S�	�s=^�p*�ء�"u0��a��}�L
�$���I�S���T�1wՖ�@���cHgƐu��p�h�9�K�WY8�q�������k��1O�M��`Йh��b���B��Q��[�}/_������}���}>���(/����kp�pcS%�Z�3umл=d)Խh��b8X��@�۷�"?X���O�&�% N���	Wb�Q�WD��/�B?J���v�cw�v�('�P�l��#��=��9F�')�2��K�q}&*lE�];��K,q�K�d?��F�z�Z�z-5��֠F��j������h$!WPc�Q>㟭z�f�[�~�����ef�ט��"������m�nl������7c�}D��玥�a�t�3��ё��KBg<T�(�~HJ�jϢI��İB�^��>����$����ϳ�w���w�����x������l�R��a?��&�σ?ۙ��b��4<����y�a�;�o������?b�I�d��	k�{���+iDD7����h�W7ko�.������zi=K�ig؍:'�|�˻����&z�o{��uOh��27�zRw�!�g�}���R���G���*<��m��{!�P�ޓTX��,�7�I3�!�|�U�<z6fø>��ӽ��+i"�C2u�5}������K��K-�]޴�B�ә������ہ�I4j��W`ʯ�� /�`s���\�?�/Y��2Tz�'��+n��Vs̈́�4� X��-�g�n��X3�|���{�V�����x:�[/o~z��T�բ�	��-丂���a�=#�o^��J�t&�C�ϼ�O�Z/�o�VJ�֞��.<���(�䢍��ztH�0�Vg�R�9��[%�`7*�PJ�{���Ql�e�ٙ���qr'B8�����Դ�]_������O��,Q�N��f�Qf[țu��^�A���~(�����ýC�����V{O����$���whI���fC�ozA���7L<!u1@���9o�����7-����dg-(�z�2�0c�%-�1a�9P�*'l�ϒ�>�r��IOx���VJ5]� ���-7��]z�;�ɺ=��{˶��
�b
��hW���Uլj=�ի:U�����NRt��~A��z���ϪF��>~.��fu)��7E�un��+��v��y�c�}C����vs*~����Ҟ��:�l�O��C:
ΐ���p�	�ߠa�=�������tх����	'\�A��]�������=�(I�-.��]7pȷ� ,���xS�X��2��I$�e����9L`T��R����Y�Lo�dC�`��L�tڛwmlj��W��S}�hA��G�[a�� V�8��	_�U�~�Ŝv�]�5�F`uB� kN�D��@dF��D��7Z��_ln�):J1uYd:����a���}����0�(b]�@�H��~/����2j}����G��Y�VLB�!�e��U��=_�������kyک=,  ־7}��� ���
�MOK���6���E���������r|~��W|]�J#@���>2A�lK�1���gc˰�G���퉮�&t� -�[C��}�����{�m(�4fK����Z��ob���|�r_!�ʠb�J]�-�35�7��6�`G$]��������"T>|:{C��N-W�E�$�=�����kO�#"�� z;شV�`��a WSF ^yI����{6J>�2��Z%��� ��eZ"�J��xD�?O7�d�g�Xo��N�җ;�K/�<̰�ͺ1���&ҟ�(�,��k�^��^B���:�������4��`�n�ڶ\|- ���U�E!�˝]�C4�Z,�����H�U������k�oQ
ؖ1��V���X"sE�I���2���̫�!��Oc�~�������~Bs�!������W_�b�K<c��g�⸫�M�ˌ��g��������϶�;���~.p4IN���B��F
�:�oO�ބ��S��k�,3�t��JD�D�W��m����������S�X��ϲ����:���]{ǷI����Z���:�����u�|p�Goرd����i=@e��7�}]�8!*�>0�~�l񞹹���|ʩIӠ�whQ"~��(�&$�:�A� S]�y78\�蒾��-y�k�>�oC�[gƃ��o
�p��MC!�s�?#5ހ\�fV"7��Yυ�Ȯxg���Ӏ����,j�zs���tԻ�	�\��S�F)SsR�M�F��'���;����D��"!��<����r�i]�	�M���M�[eJ�Ž�0��P"/B�z5ڎ��8(k�j�����38���}�}�}����N��&� � �Q9�$K mh�0z'A���\�W)
�p��{�|h�>j�����&F`��U?V�G6ͯ"�{�]��,���u2Z�tv���w�f�W�X�Y�RcCBX@k��A�?bߟ��Mi��B�)�eQM8UD�I�8 �2���
�P�����R�n��ۡ,��ȁK�,! �	�O���Hk�5!���T1�ϡC4kZMߎ��4����H22��ƅϕ����89>���п7Vğ��Y0+��[ˁ(>�o~�g]X4����5.�|��[��m�v����?�Tus�S�}]�""�{��)�XrK�,����V�,�fr�?���A��\��ߔ��w��h�j�6��|�f��,��<he��ʡ�������g@4�6_�s7��O��'���T�pٷ���k	yu?�:$�+��H�;�62<kd��٠�y6���-�5��0�<�U|+z�|?�j����"��9M��%�����*�#-�	$W���eM[#�������$+7�nc�T�Z!S�%p��9d8���^k��ULv�L��L݋%�`�����[��'\��%����>"]%nt�!9J��Kj[�4�1Б���0f��Ƙ�_L0�}h)%7�_M�$�@c�7�`�M�,���-?�1>�''�:�<vDc���!�z�I=KWb&l+:v�!��0Dl*�(��@~�ֆ� x��I��%����� �'��Ϭ�ۥ�L��@�!�Ɖپ>�<���ì�eg1�u,DS�/H�Xm��(~��o�3�lI���rD����;���׈�9�+�I�Q���쇢�F+)��ݝS�� ��[��vB*��>P^q�ܑ�ED�[��b��	]ssj�P��_I-���ʁB~�g��R�Y�����u�B�M��`0��"o�)��r� �#x>�Ny��#�g|�,�1����D�p�ɶp�sX��sЍ�j��i%H�|7�=YE�wu%R�z�c
�Ig�7�1����6@Z�����I%�Stay�'C�9�����-�o�h��:��z�X萜�X4SF͈,:/ ��Mґ�B`[%~�6���k���瓎��| ҏ�}/��Lѥr�4gŲd=�;
�� ��t@n4lr3Uv|�;:�P�,���j�/\ۍ�Y_)/���_��\��>�;d��+ѓW�#w>�3��ƭȟZ��D�7I�F��A�:KGֹp8X������Mn�@��O5@�.~��A#���q-���S�{�rӦ?c#*$r',�q7<��Vc7�g'6�[���4�-\��M�����K�-�q����а}�<��	�'��3gR$�=���Mz4>��'GIu$ז��}'���Ё����	�`��$��l�he��
?/0�SIn��{��0-a��>z<��TU��,�� F���Hi-���1w�PGuᘏa��W�[�T�yŴ�Vc��^����O���s��t�:ɅЅ�d� ��	7��r$��"���D�;����q
'�G�[�IsMc���c��>���H)�x�0�د�� S�61�ײ��,$�mt�Uբ��m]�Q�$Xեꘟ:5�b�o.�O�0x�g�c�4���Y��k9�&�s��ST�7\�S�mXR��W��VHJ�:�4_|� ~qWN�4�Z�E,#��M��]�y������O��2�<��W#)	��D���V �=(YG�������f�7���@
/��
�"�R^v���������p����Ek���/=G$���e������B�EHF8!��^���/���4d_�G����7���xD'�dޚ����3	� r�$�}�%�S����=RG�:s`�������>��qm������Jf�N�w[�*��)nD���J<$�MW2i0��oE�ٖ��UNA\��>����ٷ��Bn���jF²��n&Z)��?���P��ou~JF���}a�hqCD+�"���98�*�<P l��3�$���1�x����������I��mQ��~;�ؠ��oЭm�@����T��4�N���L���Qم!�t�#[w1�2�g|<�GA����[�Xg ��f�|e�oދ�J���@���$��Ll8M��y��*�Aq2@:95�/v���:�SF��<g�=�h���y��z#�Bȝ���;��Yb���4�#�����h����C0t�qmb ��W��/E���t��}���ȁ���22�\f�$*���No۟Џ�lYk�ډ��٧�@���"h_u��Gt��Pu���(�ܸG�J:���^�c��L�"�RP�� ��}�kr}N��&b�����H4&�fp�7f��W��3?%� �?�g�ģdO�v
̗�4���2Qf�q��b�E����S]x����A�d�<R���%�/��d_���B��N8�׳u�ȋR I�x>ɣ�ԗ)���d �5����f�2�Sxtp�^������]��K�ᢴ����(@�i��}��>&�$-��Vx���<�����8lA_Ζ}�m5���L#��/�֧ދ���P�p��xc�pQw�Y��P���iD��q<��
+��o�1���$��`0^��T�~x? R�H�#f̽�l
!�B��7o�J�0��_����.ܸ",C��N�>A5dߏ�>5��o	^o�D�MC�L3�;��5�����k�O����V\��<
��0*\�b����뜝��.[m,N�GD8
؍���:�D�<G��滜1[�߂���{`)&��t ��L=*
�X�w��00U���@�]�c��e`>(�͕����X�7��Ùz-�D����w0{�fw:C�X���6����LW&~�4��xod|�]ĳ�k�b��U`���il��KV�
0.�<(g�$a�u�%�C�w��9-�*���2���6���Pg.n����=���1��3l^�EUt�#|3�V�Z��!�QF�Laۺ��eU��K�~�q%^�wf��ݾ8��ia͊Ծ��4d#d3�oSZ</yW�d=�^uY��F��G��Z�cKa&�I~s���!$ݧ�yy�n��ع�ET˿+MK%.KE��noH�:"�J���*��j�����JT���>�8�« ��_Qn��G]�,g��騲�\�	|0�n;���j���{�A���lTZ䈓�R�ʯK�������d7��P��=
 'XRrf'��jե0ig�����כW�|+袒����}�����샽�,ET[���iH�F�C���"�f���K������vt�=M+Ykf��y���P^�Bd�و��r�#����<����&�Z�����ẖ���n�ۑ��W]�p$�	��|Ʀ�$����#U�/�1���-�'��c}x����+-���n���C+������Z�3a7&��oY��^�<�!a�}��������	萐V�D�hRv�Y?�����4��1(�Hvf3���?c�u`p��˥��x<�+'Q�]�IF:ȳYy*�G�"�壼l������l�il���B��f����w�M�-�~����(_�e(�G	D����Z�Ǹ�W��ճ�Oe�e��=�K����IQIn	z��&�ĥ^��><j['��|͛�s%N(�?��ё!|�Wy�3��9v;�i-��Te�HK���������rS1	�FL砋Ώ���
�Z2e�滅�U��Œ�&
��R�Z�.���h��!j�x�aWEf�ߦ�,�D	�2Ă�T��&"��lpi��f�-�><�.'��?������*c2"#�X�w��r����
�	��j�Hbl�>�Z��m�.k��Y�U�濈ي0��ͅ���'�þ{�BS���^��v}l2?��`��BKv����;V�(�n?)k��)'���e��j��Ʋ���=眠?ӗ�@�Fu�g���uGoB���q1�����{NX��T��}�u�92d��t����V�[W�7gZ݈y���c�}�E��R��#���C+ �/�/���=�*�/�H}K�q���.�1<D����z�������y��U�eP�+�F�R>9��׵%�Iz� ��T)�9���d1/��i{��बt\����ݥ!]t��ڍ(���J×Y�6��
t+q���ݴ�Eu�ؘ\졕����%�ۅ���꣍!��O�f�}ug0	+=g����6Z��^����$jhc�թՆ��%-�"g<��gΜ0�����"S�Kw����n���e�y툀)߭����?䓊�s��ɩ�[#5Ġ ;^7e I�Ԇ�?G� �Z�u_�R���9�y`�l����H��OJ�}�;D�V�����LAs6KO�����F�ݹ"wy����,f��JJ���{yKq�P:i= %��d��XXy�㿏)D�� �m�e��3w�m>�b��-���q�/zz�9Hmi�P����
)�9+����w��?b��8[�?e=�C�qʷAa����������bw{��vxϣ���,H�|���'�����Ů&P���
�9��'��tXK�=2K�ݰֵ���Jè��I���7�|�H: A�-MTѯg3]p����10�ؖ��^����rie_ر���K�`|#�k�]p�n����+'�����Y~Y�@��g�;����#Vi�^�ք��y��z�U h.g@5#�kiUƛ��hkA�S�c�� )av���MC��v�$�Dx�A���h�F��#ݤ�����P�@�99�:��k"j������|�����p-�R���:�M���R!A��Y�ܒ�_"/�4�T;�������k7����O6M���~����[Y��& ���ļ�5��H$0�\se����/`3���h�ʘo��!~$HU�~0i����dr���r��I�#���O.*Ÿ��PtQoD~�:D߼i����\��(9�	��:bf�X����P��OF�&j>=^��Vְ҄<���Hս��*�R�!�8�6��*�!$���h�;W�{�jl�r���+KǞܭ�<�zC�Mkia�j~D�]H��eZ�Y�եg��G�)�c���!Ve�c䌇,�{FzqY���+���5!��T����%�j����zR21��T%$j��w�vA��c�&�3�t�G\=��.�T@o4Y��C{9�`mR�[�r$ 5�(
rׂ�\��N�t��I�_Ol����"������n[�B4{��G�`#��j�_�j��#���J%�4^��G뀸x�^���`�������lH������O�A���z�yz��
Ƥ�)��x8��8=Poz�I���Ά�M��^D��e�Pܦ��yD���yD�<uL�0z���ٵ�킛h�|!`�@�6a&�^)~A�Y���0A��T��0׶{3G�81V)Ĝ��+ꉗ~�h�h}\��#Z>6e�9�%����~��s1���`���B���1���ޜ���6�v���G	"e֨�b�����[Pѱ���!���������T b��x�_z4��`{��&.(o��w��:����jzW��#����/��#�nQi3Z}��׋��.(�c&A/�r3�\L���s�5��&�2}.*8"o~�3��Vh0 ��JT�^�/�k@�8 t�*�3���YE$0,U�S*����+>�du��?���t�t}ay�=%Í3 y�%?�83��:G�!ć�cM���U�[W����q?����A ��ttE�EYv�����K3��9�/V���
y�˭�%�"�f��iKՂ�O��#�m؎S�d��wMU��7c�v7��� �aMs|�-��Պ���X(op~�%ϱ�(.����)|��$Z��E��r'Ad�����CP���E�9��Y�p��:a�3OR�=�z�Vrۗ�v��28�
GL[C�"cА'. �E��w=�t��0N׎g~�mǍ�FU�U�6ȳ&�G`~��d{;�y
��j`�L_r�:�!���l�R{��4�Yˤ&�:�R�N� ��Q��83>\KFo�ZO�-��r�W��/����T�;&�.7B���y�n7h�iN����Eߥ��X&���!:K��a� [�Y�nQ$��}4aĭ���MH�-uNi�P��'��󠮔����H�Q�K-<�	p$8�$H1�.�X �Z)�U6���H�Z����#��Ђ��G�:Ki�����([>���{���5�8����#�lr�P��I���(˓���D���DO5���p���������;O*&��~2ŝ�&�B����tVȩ��|?ؘ�0����.���o9-Im�Ϋew��{a�.�����y�fh�{�W=� �l�jv1,R�4����9*=9ɛc�OճfW>a�2�%�m�=�;;���a~�L���>3Bc��	{��;o�_�c�u���]�sF�S��N�'��z;<�m�&*�_l�&>��6����H`iw'�e8A���ߛU5z�puvXs"9�����t���1�>�E�:A�(&�e{��V�T�����F6ޡ�o�M)���G��3?1��y���x��54�.]�Etv�=�ؐ��%!*k3�vK�2�7���k�]�ܠC��Yd�EH�0�����C_Cˁ�<i���G{)Z�斈�̶N�ʤ=�&N�*	�Nt�nj��_
{*��V���v�ĬZ��uR�r����Zu9�j���Z@���������ځ_�`}̴He��y]�ڸ��6e
RA�*�HT�6��u߉Z3���W��\�T@)�UȾ�a����Sδq%n=����C#���J���QR��.a�!������8
)�~rr
TԍATl=���YC�����U�#��	�H����A�P�bه�c�V�Z�E��p+	�<]��Q�jי.W�0������iԃ���:�{]'�nO� ��/L}-�;J^ܘ.��������#-��~�%�x�/���̬�TC^���5��1G\��h�P������N�2&0�� �&�M;�P��gp\��T%o���$��$\Ǹ�:!#�
ڼP?=\��.�������Бc���̥�C"��SG�t�6Z�#u�O��T�fj�o��lF�5�c�#6�T�0]#-t�scxۙt~%������Z�ӵ�cV}�U�4���_����T��ES	]�I'4a4�O<��<�=�5����} a�@������Nz�䉨�祁��:�:��	��7��W���ߪu�F)[G�y�`��ā�ؼd��Pc�����x~��I�������P���"т���s��cc4&D���=�h�`-60�K�3(�A�v�7����J�e��)�ø����#I5�'�e�N����:�^dg��Z4]J�T�';�B_�4l�Ĉ��geכ��>�Ѓ]0r��=V���jy�(�V�q)H���'cX6�>N���'I�)��l�h8��M3�B�(/3�:�f��M����H9��Q\�︹�ډ7V�Z7YK3)�5���
�f:��O���,j�):[>�]7Ze�F�ȩ�`���l�.�c�6�E�dKqѹ��[��T�C5i�h|rf�_]�P�t[�"7�J�#����������D�+���Hд������P��C2y��s V��\��H�� ����х	��H��M5/X��9ǚ������&�
Բ�	��݉Ȩp`��ý��4��O�T皦w���j�)�PZOe��՚@���e�YB|�aO��5�>P���3N�K�]�&�Jj�\�!%��0
נO[�i��)	�W�kw;JfRi_
[�b�~<���������αƿm����3�̉����c� ������Q�I\��ȏ��q]@�!����7I��km˹�
���fR*H��r�Y��q� ^@�=ٿb�
h�����=�z .��u��� ���/?ϱI��ǩ���#����V�Q�T]-��$�ͱ�1�_j#���6T�-R"�?p���j��������y��-	�ς2�xگ�tb�$%_�|�o��l����Wk���[���(<�!�o���1 ���k�U#Z�̞����Y����6��ǐ�
�=��,K,��H>$g7��YJ����<":��z�kCf�5Q�1;Yp���>B�N��`	���55�z��DZ�rW�7���Ee��Y������ �Qj��B��M_ZԨ��pY~-~!�G��N��ꠊH�I��e���mi��H���T�/onꍳ�UmR��$e��u{�"����C�x�3�A���2I�����@.��s���,8�:l����\�С|��0���Aݿ��A�o��E3P�r�E(c^2�"�kf
���.x�M0�U�'X�l:�Oy�:P@g] ��WK�F���3's��Z8��kZ���ǘ#5�'V����G�}�D�����(�i|�!����M�?;�8�+}$eF���?a��'ï��ꪯj��-jQ%�\�h������e�yA���w`Lhh\��N褓QĆ�y�7�u��p���`gu�"��p|��7�u,�=���f�gȳ�W�go��������̵֟ް8~�������+�4bP"�lI�ծ�b,sZ�������'��W��p[�B�q0~�@H��	h��0������p��f��	c���#�q%qS�§�Vׅ(��S�]&�k�M�金\��B4�����d'�M#rt:(��=�����>�$�{�L�� ���L%7}��GxA0���3�D��� \VB9F�~������%r���ټ1X�_���jA֏��h,�shτ>�ݧW�� �׫���3�p����Kߌ� ֎��h������`�89�C|��P�g�-�K�PU�� g�~c��펍�µP�8kCͪ���-2�����n�9TW����*��)h�:�Cz'X&=���cu,���:���I1mD��I�(3`,�o�<�,�~(E��f�zq!-�#X�׏"jt�y��%&&��o��vG	��j(�s$����6Jw���+�)'pڥ� ye��~j�9W\�����e4���\Q��ʄ���+U�+�N���mzd]r���� �<��+xSC�Y�`���G� a�;�x�޶��������0	�p�͔L�����`��6a��ǲ��z�� HU8C��S�����Y��s'HX�T�~�>�	�}gF�S���΂ET��`@C����[V(�ӵg��jm�{"�kF�0h2owE� Z������yR;0�cq�� ����@��w��뀦}��H�B�A�O߬T�3`���/T�gѥ��/!*�/ɥI�hV��� ��x/���i>Xh� �L�/V�s�\��_��0��V
RK�F��LN��ߖtO�Q��9�;$P��Un�01��&�F����w��v�N���U����7�c�.��62HM�=�X��&/�C8Ie�{LP`\Dkζ��FRS��<�nL_�˥�����B�7�7�l��.	�ck���-7������a)���ov:楽<Pj�KB���?�i�c�ɦiJ�n^��� �g�����ö�782�9�;nt�`��ٝ�p	�y�F>��A(�V'��T
��yq�"� z7\?0����;w�ِI��M%?J��$�5P;����A`PM�^ϔ��C�Cw��4xA�S,/��~�}�i��g�E>� ϻW��[h���0�Da��aA�sUo^BҴ(���B߭��|ƫ.g�������)8�WQ<��;�y� �)�ך����� Ư07�g�դ|XH&�퀊�Ɍ��|��Z�&�5�c�z��RL �R�#����|�����ӫ!L�UԒ��r��@I	f�՘'�gyn�M�� ���KWVx���B�f"�X�FPR�VF��I>6�Ӹ�~w�R�C�$����Br\bA�����oT�&�2Yn_�1��!�q+A8o�s�hZ����%"�������a��K:�̜A.��өĦ�+	�o���b38�D��]��U�) ��#a��JK&&�����U��I��U�E3
wv�W�;����2���n<���i� $H�!�ӡ`��$���K���GO8�ӡ\�������p0���%�����JSj(C��B=�\���YJΆ�����0̹x�wX���gkH�!��ͥF/�H�86��"&�b=!(|�y�nP�a��sC�J�wTC�H���v�{�KK�QWd��U���������C��}yW��?��e\ *�t���A�n�~�6}���/�Α���ǺfhI��,Q���o����Lu
t�;	C�Vw1�BQ���dH����ޏ�N׿����j\��z6=U��e~�#/�f�*�[��r�8u,g[�?ƙw�eWڑv�e�)���~wG�h�-�ɰ�lXU�p$I�a+�v�Ƿ&i��� ��Z�|m��Ӗ�"y���Am�"���%}�=R����s�-������!-�@��Ͳ^��^.J��ν|�h���NP)/��9�s[u��7�0�=-`k�*�&��&�bs)?���^C�Q��A� �
�����n|:�xזvy=��h���M�� �o��|;�ǄH�2l�z��a ڏx^��#)]4��qW��g"��*diq�=�r��Z�����֧S90,~�Q����N�0��+%(I�E���;}I��A�HĐ�/B�j5����$&E��cW��LoxQ��v��F�ai�&�F9��2���5���0yqCwb�1$�K*Q��v�l%'�鶕=y�-a�oD�QE�( d�#*�j6l y��w]��,�!lL}�<s7��fD�9S��z��&��v����yKy�DR���^|�i���y��g�W�G3�^H<|m�C��x������w����07��������q\'Y��[�}#�&+�Cc���`S]�Q#����EZ�	)�Fr0G����භe� -��7���kJZ0�	»\PQ[�mH�������r�$��fn�o��=�u��njV���4�'�c�f7B .�}<A�3@�x�JP_I1��>�b��_��̰�	�@�ݎ'�I�U�ʽ��9�)(�J�!����-�{V���[����"!�q+X������T��j�c�%<��Lq�~&Ⱥ �Ni�H�r�G�P:%F��6sC.&p��y���	,����,�S4�m�Q�n`�K6��lr��VX���4�Q�h?nWWD�L%�;4RO��>�؉0MUã����߇I�6(�uǁ	�K��D�'3��56�!��?%�%m�j{Y��I��Qq�ua�3�/Ι�jjح\�ֺxӓ�M(��i�ޤ�b�kIj���z"��p�Y܈�C��]L�Y�,��A����҄^�:�f�����q� �Uʹ�n�/��N�"�Ye�T�+E�����"!�܆����n)B�*�V���|�Y�YS����f��%rz'~�}^��aY5*t�S>�u����i��@�&y��F�x�<�������-������H�=��Ǖ�5{~0�[�����ܰ����a+�+&2"¸�m�>t��q�C�qF�#��'��ɣS�5��:-�w£�\VեI�}(��#���u!�82M�C��)�o�<32!�L���g���uƪ��%9.�����S�,��ڍ^0U�eeW!�~0&�}�zl�_P"��[ߎ�{u9.��wŘ�6 ��>˷r�e�|>5�lw<YT��.����ї;O��
i0����	h Ż�Y&� � jD�Y^�u"AG�X����ug��g�3���L�_�G�I^(sy:��f���NL�;edxDn�YdI"�j���e³h	�W��55l5Ϊn-ص��脫�M��ymV��fjkU;�9�m��J�q���uE	�ְ�}��$ҌI��q������<�{'5����
 (��(+j,uޢ-2i#I[2!�au%�ӟL(��|
+�[۴�{��x�Adu�ڬ�3�|��D�O.�y7c|�o��fr��?@��/�0��&�*��
����t�M��:��xs��M{F?�Q6�o�s���,����Y��`�}FVn�1-�ikv���:�Ϙ�0>t�A�@3�.�̊����O�)(t[���?�8���(�T��'�UPY�����%6c[h>\�M����|A���(	�s!��yA0�m!eGBy(r�<1�@G����H�H��N�=�ϐ�Q�ir2Z�2��W�O�l]δo�)��q}�ݣ��A�.jaa�c2�cd��s�_�++6m�06V�,����*;i䝦8�O^�U Z{�&Kʓv���kS���z�\���4���0bD|Ad3�"(Z���@#�qT�:�
��G�c��%;��k*OX��?�C�G�n|�.M���`-+�)�@����ȯ����l�R��SH�M�_۶|6~�R�Ґ��r�{u(��cO����N��d��#x��R�ׅ��/@s�ȌK��Ț޺��(֯ʃ"lۙ�	��M�P払�,A����;�f������d.C���5�>	��f�<���y���[N����K�z�%}���U��{t;��C؈Rl����hPG�A��`
��Ѐ5�C�H�|��g�?i��ۢ�Lw˪�2p�X��R,qd�����*�(W��FB�Z$���eB݌mq�MWq���*;��� t!"����9��G���N��_��z<Hw���S��{�.-~�2Ө�v�H��+�n��wNji>������A����F�x�>js F_S�1���O;cNV~���(2��" Ud�:ϛ��̌!J�t)����!Ӟ���9/u�@���Q�������Oc��a��5�R0rzڈ�O���b�}~��J$�S�~"F��xk�����9�3����>�B��5��*[��	:qJe��>wm���r/���6?'���l�n�2&6�V�:�-C�5�V�#V����U��}��/��sΖ��4|B=��UbY�z��	��^B�Hnr`)e�:XC.ސUB���F�,Cϯ5~���������z\���.��܉��p�@�A���26�].�e�ƂJ-��Cڢ��W��AR=��7sv='�^�%�`h�M�k/�LQ�g~Κ�{E�A3.����I��\K=S�mC���m�f+��LRV;����ud%ߜ�^�+���7Y��f>h�ʺo ��'4�g2O���2=�q�U;�n�R*���%��Mb��QOv=�	À�Ɖ><J,�Rn���}�]a!c��ן����A��<7�����Aު"��x^��[H(��,e��T���KJ�UxA����ARv|���E�?���}�`T��b/�H��	t���qG6f�M��k�UU���-���R��"�^��;]���Y��j@��Q>�b\GZ�,�UH-?|��<�L$6�G�tǘ�$�w�}u�]x��-�$�# ��--�B�c4�6^�_���������|q�De�p����S�g/H��� Uꖾv��ۻ�p�p�'�h�?`b��`+����O�4�1؆ms���O��X��D��x9\�0�24p¬��m�U��lx_�8,+x����}B������z�X���V��a㽴ڰ�X��`�v�llbٙ���Sh5�����މ�;M�<�r�� �i��_��#�I�sB�LNS�H��&���=��-Ud���n�����?KCv�w��{nq�rrT��@��6@�;S���xL���_}'���������%>;Q3��;�"�C.}࿉�3������9�`8��e�aF~�2�����������-̘V��ݽ0���y(���]��(����<L,ŤS����M�U��hg<�8�湏n�Q�6b)��Z>���鮝*��$�ׅsKT]�5��7{�A ���Ij�՞$��PL���D�j�D�lX��	���w)��=��z���)�Z�Z]�������[J�X��>ި�1��<�ߜ�m\v8�;��� LE�I7q4+���;A�\���6=�]m�V��**��I1���������&He@
ݛ~!�ű:_#aU]ѭV�/I͏,}њ s��܉���I����梫*v� ����&��V����mi����0��|� ���'9
\S�am��'�6�Do���͞H������X* ��I�vp�[��=�$T�z"�e�����Y��t�?���Rbo�E����[֜�,o=�_蜥�X���i��,/���{|a�Q��։h��
LA�ߍ���}G�PS�����~��&5�7a�y�"uArj��2�<�5�>)6"M';����1٘R��cl,�I�(�z���l���L�3���Lq*7�=<q��G�d�o*�������i�b��tl�
f��1`�T2@����Is���
ș[}D�"�Pr�1V�KE�9 *�]��a5NꝮ���8.�����2��<�+�nͽ�s#�##\�p_��v�к����L��@���X�r�
?c���螸%�!y�a�^�cv���M;������9�TJG���U_

��*��+e�����!���0��"";yYy´i2c�t,!�^�tb����=3��a���I ��8r(��7Ȋ��H���o�pN)RN�����t�|�K4�"Ոy��͗KJV��$�1�L�"�7��r$��5J@j���
����h��TIΊ7 �~�=��?�������n6�ҫ��=?f���#�]��̗��2S�o��5�
E0�mtj���ED66��y,c=O���j�G�v��FN�s|���
7mU��f[����34�l1�p*���홷#3Љ�{� �?w ]��S��|ޮu]��h���Y�B�2;-��M�"�_1��҅QN<萪m����
�t^����WW%ЭxnW�?.��� E72�%Xmd���{U�E�|vrf�.`��~���bya�栋����S9����GnMv%~Ѩ�b\q�9��?�>AS����?���f(m�B�S�(�*��N�ݶ.�����'J�,���t>/F�D�ɛA�{y����Up
p�
��?;�&�����V�]�6��/��]����{7�+H��^���J�3��nW���!ފ�r�H� L@���A�6/)��W��ᙘ�L� �$MY�҄��
:���tT���gS%��3N|���ЛFZf�$�&'Ѵg�D_8<���M��z�p��Vj��$Sn��?a{�I��<�م����y"�69��R�����y5~=���m��wT�]�>NZ�sq\I�](�����(�(j��Ⴏa�9g�������埛�*�'�|�z���u��͏ъ���d�������W)Ԭ�_�n,�P�y�Y��b-�}S�5p���_WB�6m��X���=�T�)��Ǝ���uS�K(2�!��Y���L�G;�h|��,4|�JRU^��去���ccRmQT�D��Xe��-��:"��'����D�O�F�R ]�c�ޚ�8 ���岫�rY�}�q2��ph�@䑯�z�v̌V�eY� �|�����ߌ�n�G�d�����L�s�%���~A���S�^��|�����]�An�Aubߔ@V���R��5"���C���eun@��XzSji�&���K���v��+��4�1�WT��z���b����k���ʂ�x�؝b��s��>�`��=�Fi6�/5�KQ�IQ��^�I���>�C-�u�ƶ`��>L`������_�J]��p����E�H�)n�Q3
�9=j����O��q����-�ڦ�)����g�G��;^���3��,��]�.���7��$���W����lFӗ}�{�n.���K�}a��3�!�O���d�{퀸�&��� ��ag@oD�td�GE��PR���K�\%��.8bX�,᷍j��ݶ]8��k�y_R���`]�|��-�Hg��M�>��ˠ�eV4Xܵ�Q��إ��/���s�����ö����M^O
,=>0����+�-��{ J�%��p�eǮ5*�B2�������V���c��'�Hr�b�6>t��ϸfb2�mD픫��s�b��\(#7JX�����_iB���0ZR5X�ry����-��I&b�=���$+�F&3<@ݳ0s!��9����F��n0�跙8-���~��os���9�Hw����$ˎm���F�� �@���hd[��H�CiǬ�O�uS`�"1�`t"pʩ�"k��v�J(O�WC5�1�q0ͭ.��DI�)�@*#���p/H]�m��Kj�:tԍ����x-%�Rc���s��0���K]bA.}�Ò���b����ܩB�E����D~�(|���9	Q་�n�����g�gx��I+�Q(���a3W�� ohZDcFQĻK~�cਸ�Z��_c�񐞛�?�;#q��k�^�fK�Z�ǯ�T�{�;�vq�-�e���h������w�؞ɯ�&��p�r/`�xTt~�T�dpBGX��NU>��OG��a1N}I�����򰪜b��b	��N����B�Z��ܯ갑��k����0�/�m��#�T��U�w�/t��	�䳿!}�QI�H����������KYnYÍ���榽]̋�Е����e]�/O��Ծ�ST�e�K̨_��I/˿�)(��y���s2^�9Z�?0,<6�2y�����5#�6��t��r7��E����E7[�y&B�j�ߒ>\웷����"Y%l�����e��0�5��� �E��or:ɉ�e��-!{��2�B�<^N��������c :8ݸ�x���0v�Z՜���2�e��ZB�x�� �{�����iŗHn�H��}[���B�P���0�8��1O�d�g�8��U��>�=���T���p;����s�о�u�갯�G�j�2{�~i����d܎�{��Y|K�@s����<X�5�oO��=��Bp���6'F�R��J�3{��*d��B��m��:�<|�-��d��)B��ٿTޣ(\����=O�֬��DRY�[/[��B���Ü
�g`-qu�8j^a3�Xݵ-7��1��|�~�Y�!Z��>v�$�b�㍃�ZY.�N�h�4��(v���KWIX}Z��t`�A�qe6l3n�3$�?����Q�)���K*�U�Oo�7w��ّ̏#�~6�q��J�Tp~6T��̭Y�@�Dk4;���&��u���]�c'qlhҪ��%�̙H(Q36gP�=��m��\�3��������3m=32�Ƹn(�n�vM�:��3���m;�Ӭ���ڷ]c�j�w�`�o�ؤ��6�Պ��.�M�nΙ�W�+��A�i12%�J!�>TxY=��{͓l�_����7���bFv�0��ӫ�1E�D�w�w�+,�ª��8�
ol��y"� _��f���̇"ղDP���bM@�i�W���^�܆1=��iA*	�@x�#���H�%tr�|쐰��B2P����ܾ#M�����\J�Q���2�5\?���S��cc/x�Tf/jN�����\���gR�o��ڸ���-�����m���t��량}C�z@��+�����0�	���N��@+�21�����}�N �r���F����z��9�M�1)�A�-���VB�m�T����UB@�_����\O0�K3{D�w��Om���Gm�ţ�
I��R�M.�l����|��H$��{R���M쏍W![���	T��6\��j��ҋ�[;jJ/�/�܏B��;U��1c�ll�K3� ꏻ
���,����ye�潓�lɻ=��}'*���er���n`��p�G7AE1=?>0ѽd���Fz?,�f��7�ph�1�)�Igv�x��j�/���[)�<$�CD�n0��0�t��lq�	`Չ��'*�*�g���x������nd%R�'&3{(���Y����@\���6�	��J�pL�FVX{����s���ra�܌�ĝ|��T���
VIҊ��@k'?U�>�G�=>fT�����+�%��x���Òм�v���OV�#�;��͠���oM��.�4�T���0��2�C�lL��V
��}!NQ�:��d�?b�H\`�v�W��䍞4K������iJu���l+�W T�sw���}�	��P�xG��Y�^��G�s6��P����	=�_���5)(����	S�g��q�S���c��� �}��V���{����I��E�{�x�A��:Q��fg��d^F�=Fa����$�}�R]��(��7&�;Kگ���Z,*7�5Qt�!�o��7�d�b��v��W���g��($12嗪�a��WtgY��jMjSg#u.>7ܔ�������mZ"��'�I���ֵ��|��g)V�>��D����P2�l�va�����������lI��$Kk���V�\��*f~�Xh��A�l=���e=�g�k0�A��X�e�=��$�Wr���e�LFL*��6ې�M�I�������o��x]��0B�o�� y�BL����d�2AI��S@[:�,�M �(t`�b� ��W�u:��6}�I�i(FV\�P&��mzʃQ A;����s�8�T�49�sm ��fD�qL4�K:��P�� .�����GPc���]ɖL��':0���A-�&V��ըcjR�_�!�,v�dv���nXۑK�(����/�#�����1<K'��C�E.jʤ��+B��m4���5�-��5s���56�k�S�]�RP=�Wh<�tz�/Wwz��8�_�x�	��L�gP+̼��[�6^a7p{�b���ZN7`�!� ¹�� m:�váp�Nw��u��g�8�����xx�s=55%�Q$�?�a��=�?���xlYV�y�Q��F+�?̅���E����y)���o��"���0H*l�;��}L�KP�g�6�;Ǘ��F2���f��#��GU|W��#��@2<�0;��N����D�!I�F������&� ����mI<R�����㍢�+zk��v�(D��H��?[��p�@H��C£G���"$��)P�Z��z G�Դ�a%��^�y�������Lȁ���o��)����G-uB�
��,�a8$@��{��8@Z��h%h Gh�i���A�&~�:��Uhv�"���������}dpUM��2�~��HM�v�h�U�W�>ꚧWW�~�����0��κ��<�W��K�t]cbJZ��,��W��a,�+K�Y-Υ�P!����y#�i�s�"���6a��?X^0y��~�����I5f�a��"��X�)���̶k+�*v]�Ю�m+�Ԟ�=�Np�[DG�X��w��_�L�G߅2A��mj2���è.�\�5f�nȍ���_�n��*ţ��UN��O�qj�F�����Y�a%�5�5&�{�%��萅	�_8&���2�P���ڣ�Z�L��iHSқLp���H��۴�X��d_S�~��t�ف`�zn�jdrV^gk�#\	�>7�oaV�w��sp�L�"o^ɱ �Q�x(�R��h23_��g
>�
�0$t�c��n#��c�E��|Q�︠%E��Ʈ&5�OXT�V��>�x�ę�9F�Ns?A���?WKh�C���-�� z��S
S�R�}�N\�J�^����fw8*{b Z����I'`�U���D�՘ӠRq�b^UvO�Lx� ��^gz��~�_.uZ�B�T�[���Q>�PEl@́�2Nh�4m�) �ӛ[ikb��þ��R�K�?�_M֭���q����g�ޠ ?���(��#�h�!iT�v<��24:�b��Iݙ����q�����K��`]��*^Q>���CK�Dݗ�:��
��~�z>e�7��!s�P��K��By�wx�����o���[�Ԩ&x�)��0!צ;�g;Ug���� sB�0)�aÕ�7s�$w*�8��S'�Cw�)ŹQ�S�>�q���x�a���~Т�ЋE�����������d8�J���#�deϽ�&P0AV���a��0���h��,�n(# ��T��OE���O~�ꗱx��02|C�Ce��|��8��MH@�#<ġ�����tŰy�0�K5����;u��,��8J�\?�u��养�ja�w�04��t���
c�y�������$@�J���;��~�7�0� ��C��� �u���_�?R����r�D�~pT�:�1
8M����VG_y=�<�wL��O�HM#`�@{�Ӽ�(�D|��)Q��E��7��#[��c���4MpS��k����!c3#��V"5�{
�,��a�x�	/](�{8�^tn���Y���͋��͢]���X]f�`"�(����C�):Y��q�x�+0Q�� ~�ο���s�`��P�\:��+C��O!^_S.���4�A7�v/,������m��^K�|sX�����.(7}��ԩ}8��c����������^��>e-ҕElV�<�~�;��\F�ܜ��u��y-�:0:�'u��rDU�'ǜ2R�%:E�;�V6��-Zp��'�[D�e�}�$������Q^~@k��FM�g?����@(^s�.�3>�<�{����Y��5E%^����ִ	7<�꤬o����J,��e�?��݈�<��>G)'� q�lV����%�|%�y*�y�1�b'x
.�|��In[Ү�]��/N[o�s��1)�.14CAf����{)�C���6�	�!���}�y/��)�xi_��*w�w��-�vi�'!��e\f�6ۙM�Ɋ�^�����aǡ���8��܈��F�Vv8_\%Z=tq�J8qQ	6O-۸Ik͵��y�L�߆�u��[vF�U�]�-���m��k�0Ơq[*�L�#�\�Do3s��ٓ�M`���z�q�� �����`�b)C���i�@�v�8��U��?<�|���4�l��Q����g;�!��D��ܸ4r1J����(�@v|G��Y�͓�j�w��,�(Y��oN�_�����=�&3	�ͽ�J(��g�����g6��{qS�v�����-:1p��´��b�ފA:�I̥����%��%8�a�}��:���;�Yvg �j�66]���vnǞ���1N "���-t��\�h�65��&���eKR�L�V����I��ʍ�#}��,NGȩ����3�)�>�ܴ���[��\<�$���S!�
5L�9���Bq~0��g:g����)�A��m�*y{z�'�F�{�����Y�%l;�I�f�+��"����qޞ��#��1��;�&�(.�,���p��-B^���ֺ�S1�7L�hU^G�ʅ�x�������P��o��լ��Ղ9
�W�	3j��(X���yBY"�N�	�=�m#x���e�D`�m3�K�w���.KP��՜�C@���Wk� �����|>Q����uM���� l3��H��H�?��7/�X�?�x����1�[�b�gJ�=���^��W��.��X�-��'>��j�k-����g�nB�$��)������2DQ"m���t�z14X������y@J�"m��r|
���/k:= N�*�d��4�SI�T�[� /'�P�i���G��j)�_�S�"%�� ��GW'g�ݎ�fMt*�Է�f]@W����B(���+.eB����mH{�]n!�7g�܋_���j�k����V�������C!�,E�y�1 4K�Nڷ�Y�u�7�lJ��	Fԩ�4�.f��= �뮧�<�Z`�V9ρ4��i�E����_J}BՍ��5��mg��E�R6l�,��
��$���Z���a�&��'�SĆ�ifl��F�R��!�SnX+��a�r�ń�I�7@#99У	���q]���)�Wz��Z�l��K��Q�+D�b�
(�u]��[��Y�;m.����_�j$w�I
Y�?�Z��[�]3]]J4�#��sL��������3����ͨ�#����]�ߨ&?lsb�z͌�R#A�f�`�xH�>�7z�.x�,������;�W��T����`�yb��0AJ�����c�;k���kǴB5��t���va���c �2�����	��M��[�#+�Q��� �^�V��d
U���{�(�;�F�n�K��'�s�K�MKΪ%�Ĭ���:�]<@D��澏Ԡ�ODhj��o:[t`�$g���ġb�ﲳP���짲m��n���7���H�'c�p��}�2�vq�L7��i�fT�ʁ���<��6$��DJ����*��J�.:J<���-�uL��p�'%;�Q�>��4"3�wj�K濋���D nBE�\�J�l����f�&h6�Ǉ74ɬ	�@�'s)cӂhd|���Nγ����i�5��`�L�!��9"�����bӆ7�(}���N��mI�W'P�Կ�Ag}��.������ 7�bqʤT�;Bk�,>ZW� P'{�KkU�Ҷ ��}��6�i�;�����?vX�,e��+5rA.pG�K<ׇ/�L�6�֋�"�.��f��k<�Z8�J�`w?��Dڭ)"G�ͺ�����D��nH�T l}N��lD�a���^<�i�2��Ë1I���)0�����|� ��Fl<AK 8|� ��q�K���-{�; !~N�k�C|A��](�D5�Q��"Y@����:�>�ͻt�j��������X�AB2�����"�@���#"�I��3�=��G*aeVt��eR�d�а�`�y�K��)֨���1��X��Ep��~,�j4�����g�MXv��o�B$�v��!6���&ߪE��8��+�˭B$���ًj}��w���[|�VxH��rN�����q8bI�T��7���~:��@x����[Y_;��<�ޢ���}�4�c�eG�N���X?�=��s��Z:�pa(�ܽM�X��3*��-��B����4z�ߩ3`'8r��>#�j��q� ����y/]�+|� ��[�V�gqx�����5B����/�ΘP�<��|[[*�UIPqj
u��N]�U�˿8"��g��R
z�Rӷ����q\q�6�`z�B 6�����ci�8���1��'��{y�bjf�����G&h�1��S0*����ak�f�.c!����9�+�?������UP�7�}I.�4 w��ȸ0��ܾ�ۡk�O�|���@���,\4�W�eeF����4��"����n��h|��Ư:Ρ���&I�o�\��i~��En�ز��P��@f>#��D�с1��� !���?��9C|�oP�s'�Z�I���@�@7��L�$��?��﷔���C
�9@̓M��Z�k��۰n��)���������	����o}��fN\��G���h�7��C�ozhɜe�A�.����o��q���*R��>�F����j��CRJ��(�:��鱖.D�t�� �9_T?�>��k�Ybb������~lt�+�d5vFLt����LrCy������ bO��.��`��96Q)T(;$�U@�2����f�`�}�Ez*�?�
8R�_�1챼�I�@&� 9_�� $��e���C��5��R)Ճ��+�!Ϊ*��bKi]�.6��� J� ¤��,�b7��/���3jIȫ���EN�@R5�ڐ�-3����ez��T�g�z��8�,�z�o��Px�
�B�#�~�HϨ��>I�a�pk҆��:�� �X���GMo�8g��Ƽ����G2J'qa���h�W����������]򀧠c� �ge:-]��T�+T��\(��
�������!qx���݁�o0(Wq�Y�gأ�	��q{�l�A�}�]D*`�g�h�&�Y�y��U�k�*��g.;�����H�6���C|׎�4R�}w�)t� ,X������-F0V"����c����*o�)!s�i#��T���m4Lnj�������q�a��ֳ8uf��=�9ׇ
�`�=�Ѯ���\p!�ti���!�{�zz�"@vߔa�JїM��L�h��)�	��_��	��!F�F�Z��ӄ�Ш4��/E��~Զ!NCga��+�#H0�A��k叙���xyg�9g������'���3��4��=sM�,.��	���J~�[pD�i.��}v.݌�v -�g���u��^�r�����*��ˮ�͟f.�