��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� rā�SZ )����C.��&0C]�-��[�3�-���+��պݣ�k�J�vo`�A�����f����u�X���v�=�а���]Q�Wۿ�߸�=_Q�X����j>��Zw�K��SvX��ƥ.���#�����Z�0���#7{��\S$��@1I�QX~TQ�E��db����۰� ���>0�%�9�j汈��}��1� ��2���h�G��SeY�a���	'<x�p��k�H`�H�j^y�0�s�78+���ֳ�`�R3dW��_��{p[�?$�s0��#�zS�_��bH
�c�p�IL7]� |����Q�� ��Rr���=��E즕2%�����`�^��l�q-�]�p��jf��Ӽ-f%H���ȳ�>��+���M�71��4_�) 3�46h�rb�J�W� k�h~K0�>P$�_n)���5�r�j��W�J&޴o��$>��6��ŀ�;A~<6P��K�~��f��*I
�Z��}`q���ApC��n���g���3��-�іrO�mF���,�$��@�BI�q�}��Ȥ֐����î�䂧��@������U���vU������ �T#K@f�㯁����|95<@���+�-�)�����K���FI�k���*@�m&���
���ma1[�2�u�I�\�U�yu���o�|��2����;�W�W�}P�K>%5�'�8���׫=����k��,�t�M�0�8]q3���Nܺ�^�5Xz��t�l���&��}��ޠ=���< ^�8�$�2���c�=@Y��ɤ�#Z�i���'�*G�����*��2�s�`偞�gM
��㙘&ꉽ#��:=���7�����Տ�k���i�{��I/��ha�[s���7�^��8�鏋��C�ʜe�R+!X�"H�J~�Q���ezJ��=w6�^8�Z�w�ՕZ5����P:O����K?�d�P�z7U|�D-̶���ّ��8�dӣ��ǯc�0��e^�ɒ��"����f�V�̉O��Mys����A�ň�7E�s���'�i(1@D�n�b����οN�/�����Zz7����+�O���o���VM��)��w���R;�B`ٞ؄� o�19��m@�K9:�8I�K���R��a�2>1�4���uM 7���B��(���o���������|D\oV���,��k
�ɩt�%Ȅ�vLP� ���%��L2R���2�h�MKŻ0t�Cم��Qf� Y>`o�䢠l���V�[�ƙ��Jh����7����h�2�RH��N?��#6�ߍ�%��	�2k8����%��*��׹C���t�,��~�Ҕې����M�<}~t��+����:J��&�06 �_ão��SiB?�j��w`��G'�ai.�,VE�5:�Q]��k�'l�/�K���ʂ-�#����T+"^|���y��"�ʟ�K����_-�˷ċt@C%. Q�+��̯-D�h��^�")\���ri.Y�?;)��!��u.Tb�r�؏E0���Ej"�/'���+M`;[�!���5�i���y�n���-�Ap�̿W�޴l�x���E�5~>z_�v�z/T1�������>�G��b|�v�Z��6zXi��x�j����7�PS��O�j���_�������QC�u4�]c���6��~�)x1	�-y�����)�Oc'ɦ?g��A1��4���)tVz�!eԦu�O"T��$���$�N��M�#Qâ?`��'�i�U\���	�����u K�|�о��R�t����9�j��g��P�d�@��1p�1ɪIyw0�pԢ����	j��"� �;�
x�ot�s�4"��q�*����Si�aGv��U���s9�9�O�a�Z|8��ޒ�j
X3>/k
u\�ҙҤ;�{�uD��$4c�J�l��w�|�KM7Oc8��~W2�uX��W�eHи4>B�AG %�q��K�5��D-Z���N�����ju�Sm=�A��,ua�]��א����.LiI�|at�Q����?�L���a(M�%$�GR��>�7�)K�"G�oq�,�d��j[�]GK�x���^��KfL�nS	�)���{����C��<�e��eU�K���X1K|B�o����j�ӯE��}|���@����j@�c樫���z Y�hY���#F�k�_�`U@�K�5���TG�B�y0o1��}��T*��2�]#	�77��7r��%J!�Cfp��l�pDp(ML�mH�7R�_71����[{���� �)B�o ��raZ��id�/���A��I�Vs�lb����廻ƷmN2�y�����3�-�z��Ş�������n�6�Krz��>��{kO>I-'Q�=A�Q���~[ �Wa�2_��'�窩��(f\�b,�Q@�t����Q&�f�zJa4!�oX!�)��a������_��e���
1t|�.�Z�H2c.�L�8B�޿��p���3��I�B!�(I�髀�ʽ��W"1��\z���2��0�!��H.�Ȳ
s%L/�هdX��������@[��㥯|㋅ā!h��	��H�5`H�`\�$�x!F�[���Ao�9�5:#���(���}�Y�*�!Bm?-0���6Dȼ�X=�u���l��
^&t����KC�������>�Y���A�q�������H	�� Z#08�����#�X�@ӷ�֕(v�p	P^>S(�H|iG�[ǯkK�s�Tx�@�+y(�T2x��+�5ջs}~F���\�i<���8Z$cW��ջ�B����;���H���Ki?�c>����$�H�Ck{�9^�ۋ�۲�5~�����Fv��Ї�:�;;�Q�S�[�mvL0m[��ڙ��>�\V=~���Oю��)r|�냿?�$~��sݐj�X�Y��ѦDFzq��:��y}S�'�ru����ֿ�86�����4tʵ�#sF�S&~�g:e��om1ё,�&�a
�����{P��~��,k�q�� e�\9�ނ�}���z�`�i�0�]YEI��ϧ���K� +��b��%eӐ��&��`32??*��r����c�L:V��Qy�t;Q��P�B�y�Jy9/�/q�$���Q�T�&t�Z=�a�N�-�����0�l����>>����^�жat��'�c�G�V�O�S�+ �_I�*F`!ˉ5a�u�C�h�:[�Ƌ89HY"�'�����j��B
�³0��c�t ��f*5�"
��Tg���Q�}�1a�6� ��K�
|"<�����ߩ�V�O옢��K��=�w
Vx�G�"\�8�	��t*w�k���ІꓪQ���\����
����݆��}�)�./v����N؆�(8*,<8T��%x%���Ã�m��{�{�&5������,�V���
<.@a�)�M���j4�Jl1/!S��;���);�B�5���
a���l)N}�'*&���b�0�3�3f����������9��2�i�@`mv�b�m1Ue��w�Y�N6� ��2�F�(]��f���)6�=�ƍ���k�z��\�H!��_�U�`�LKnz�<XH�E�� ��L�����>W��8�����c�k2����1z|W^�>#�V�̵��pK#��z��(l!���^�ߎ9��Ɗ�a�=�:����_"�ZSy��Y�Ҏ�h�Q�YG�!�w����4�JnJ��c���]9c�e!�1���#��ȗ���f��V�D������������L:��<}٘��\�R:(w�l���S��%퐷����(��B�<'��R�\���������EY:���~Ve�*��f�|�Q;d���3�g�#ؓ%U�7�6�bϾU�bm�"e?>1��mʭ��Ω���d��+t��:�����m�Ľ�ыY����\�P����W�_�s�`��'�a�y���nQr{f�
��$�1�c͹L��f�2�f4��ܻ��\%⪒�:@D,��6tR����Ir�s&s���y=ZS�me�9z�~�������w�]+Y�%b{r�U�q[�>�RrK �ѿs�$Q��3����Ǡ�0�P,������l�Z;5P��4�\[n7͌��V��-�LD�1e!0��b\�����"�W��eDx.�V��9��if҉�K���g��/�/�?3�nCS��M �R�a���O_��1G(Y`K�99j�%��I���m�r�Z�yw|S2�甴+�lۢ�HR<�:׍	��O�B��`~>k�E�����A��-�>��{�ٔQ�Kinfk��Ad��v�y2�����G/g4lm�r}��v�|�է;�E��
n�*O��9��k�m6tz$���2�e�,�__�m�j��$zJz���zƽ�+n��	篧����R^&nk���:����Ó��u�Z	g�1
mN~�m��SԯY��ݲ���r�2���K��O��$��(~�\�	x�AIu��Y� ��� ��P�z�Ssڅ���g�u%�|w�����:C�Gs#��d`F�=?�oj~�	 $�ڭ]F[���s'��r�X/ ʓ�H:�i��"�40�0�v�x��q�L����]�O��"ϠL�5�|d���گ.%(A"H��I�c����ye+�4H�lJa�4���RS��c��X�Ǉ��rf��/숃R��!���rh��Y����A��|�ieMR�TG㽷>@Q�A[����t�^СDMY��C�$U�杅Y��RP�/)G8���Đ���A��:w�hP#�B��,X�6*.ĩ,�%[�GtcI��g�b91�}|/�-��B�֬Xp��{�����T�n#�r^���ؗC���zU�v;���[�C���mV6x� ���e�E���8��r=���7��_uظ��K�a˰��{H�P���U_�������J���vU�7���ՙi��2��8�%8��4��u���i�ڬ�\h<i�Z��đ/�ol����N���*_�U�HK�m\��I=�OuÕqg�Ŷ7�݋�ƍX3���Fo@���!��Q&����y�������� 6�Ї0��`�ܮ����2�2�`��Y���RӾj��䦢�ZQ)���j��VW�?�`�h�#������mp�D�;^�����sj5�t2��/\�5k����#�M2�].��-^��5-َ,�tv~�v�/ɘ�9��c���J�}_�f��s_����F�]�#=|�G%������ZS.�UL�{w��&��(�c����u(�P��i�a~�P.�<��m��u=4�Ҹvj��c�F���e5�ߠcE�Y�f��_y����t؄b�o������?�We�S��-L�u~ib�����������@� '[ߵ[[�|��?�y�����"�������|4B(�{�C6��G��k̅�1�����q�͛cPܷ.w͹�?���ӻ�kx;HN�[J�Ҟ�F������zɶ�^^,=�n���}�
�'�,O���?�4-_@��U:d�k�Q�(4�ރ>�]��o-�
:���3W���
�Z���;�.G2�F-���>���81�U���.�د��J̒���Oj���!��32)��� _ �W�=�6<RAL���Vpo�Ơ{$������,���
R*6����=�¬��A�t����9�l�J�oX� 	]�%AO;�-���G�� ��|�a��P����Zo[��N��e��p�zs�(�/��aF�9C��o���B%�!�������-�HO~a9��Pp��I󹋮�[!Ir�����;�C3�TT��A�g��!jCqnp���׹�&��>���O�S�Ɂ�Y=`崴������?��Xm�Aj�_1@���c���nR�A*�A�N��.��+Wn�x�.�������Y�.?�pyMC����+!M?�<��XV�;to"q�yF��݄�;�����K���A_	����=`K\�z�����M� ժ�kz�`	�F,"�U�m �k�	���c��ܒf�
q�Ȓ��ɧx.�o��p�).-
t���oRp�q�`ʖ�T��`�D#2)��Hj�W~t�5.!�w3@����X&�����+��,U�-���lJςؿo*���0�����̀,=Xw��3$��!���)�z�Lgro���|�"_�c+�%�M!8��	'q9xY���Sn�A��'��D��GHװ���c;�1��£z�%���+��܊���3_\4�1������ePH�0�ى�cUݲ�hG�9�ur�ƾq�=�� DtJ��������&|xbKܻwÍ)�7�����R��\>�4����iu(��w�|���b2�247}7,K�L��
�<����K�'R�CQзb�SO�!�@�`~ ��vp�X?�i|O������f�O��-W�9�1��fI�e�'oQF��
�~�j�nӻ3:47:��DE���a��ύp֨�s�|^bBkA�M�X&��8���ZW�=t�R$�����/�q�xXs�`ޟjt��).x9���҃���v��a´40P݀�Ƒ��%��i��pZ�.G*	�̮̉� �G}�@���ؚ�Oҭ4��{sM���=j��թ���ҕ�����+��nUu�U�%c��s�]�DXc�|��}O�O*р�\ť�S�n2�	0#�˳���:E�5���B5��؏|�B*��Y5.�CD��vgn�8��X���#Xl�?����m|	H,-%�G���Nd-?x�Ed3��	6�E�F9
���S�B�3��N�n������PF��'ET�^ڵ����مN3��\ϱ��|6q�������Q*όPf*;�TO*��*\�"b�S�v���֣k�Y�e\������n���ǹ�j�J�y�n�U9�����BLB�[?yu�i0s����o��;�W�R�����
��A�%`����<%�����`��%,��"/���V/�m����(�������}AH˙�) q�Fc�����mB१�s7S���M��T-_�r�r,;�}7�D~2f�tFQ{�]�'�R7�GQ�������"r�4Q$_l"]�ڈ����&8#u��]��h�k��� �1��no���A��:��;�^�>�Z�s�X��+�+�Jz!�d=��/N���*����4�6(�K.�Ie����n3#�k<�"���<��N��YF���]�d���&Ħ����u�~��ܖ�w!k�њ�Pr�dd8n�X�:�L��Y��\g�@F�m�
����B�.*ޞ�V4Ф�Ļ���y���7���Ǿ�]njV�C:�������c�҅��� �?�;��x&8ɔ�e1��QZ�k�v� ���XM�!P�h�IY}����� ��3�D�M2��I��=����q�v�������}'FF�%��v��^f�M�L�
���������3C�� �Üh�n�2gY�8�.a�S���%�|ì�Ba梥��/1�2�$�-)L�<�����<a���)/���ׇ34�o8����Z�Q�'�S�r��"�4�	��z��?��
�ŷ�%�<��C\���'��O���>>d���X�3���3!��
���ŝ��xs�&T'x�*_����*�w��֢^i� ���6��,�kX���L�r�*ۢla0WI=���D�xSI����{NO,����'��}&��-����2}����W@`�)��VPk�놓;�w�3�4fWB�f�C���%��&��ɓ"�N���?��_��}���=2?�#�z��>���Z]3��7��9L��cwU-�\�i2cgZz̩�̚l��%��.�b�)��i2�P5��D\]�
 �Ly*���Ac�e�4�!�N�m�Y/��+	 �vN^�Afն�L�&g�J������5Cs�~�L�;��N��-B^�<9����첨3�Yj��-i�r�W��9ݷ5�~2�W�<8e�Y\V�����9?j�7^���r>����!>}+��d���
��MGR���5qf!er����U�xIS[�ZkҘ�XW��A�<�E|�$����Z��ˎ	^װ"�y�N�{[R@g��H*o�/�riTuǒ��%W��#��L��d6�1TD�z�R����/�(�QLAK+����EP�Gf�맲��4�e[Hb��P����E�~��c��L�RdeIP5�p��Px�хJvXh	��(��p(j��y;����d�mT����-Z�6�$-�H��&��%��K�:X��l&��(XBD-X�(�&�5J�h�/�����}b����E/��m�e�Rv�7� ��[�=X$Q��=�53�S8��=�� -��
����mJhr鍌���z.F�Y�xB�-1t����v�]��e�����U��#�����w:�Q#�r!=�;E%���0`�&��k}wTl'8�*)>���G�I�R	J�u�唑����C��j�<���]�%fD趴���^��(a����M��*E�`�=W����(Z�xj��I�+n�����(v=��V�>�&knֹ�����υY0R {Tն�����+om�;�^U)l:GĽU9�pL|�����lZ 碶g��@N�?�FU���%颴=�rQ����+K2}��s�m�ZύNmf@��at��>R_~����Z� �ӈ�~+�!�7ֆ��E���DJ0"���N$���~�Am��íc(��� o+��b��[�hLB��������$����g�	�49��In��L&2�F$�q�,�!&��]�>m���y#�-@�ܭ��;��+��[q���)O�t#l�$V���y!d5(�8�q�����ta8����k_���{Bk��}��#��{L�3,=��c���C`����ӶH4����$Om��^��M}n/�.���F��1�c�N�l��q�'�w���կݭ���߸�ͻ��C�f�"�E$�JO7	u�!r����g�N�C�yb�O��rI�����Ӂ}S�ڲ2PWWAr�C~������m}�ǅ���nl��M��r!AK+pU�#9��ĳ!_�|�� �|�o��Bf[b>KR����>�&S���q3��nnoޅIw9x�ka}3�e���,p�G
�mkc��.p�%�9X�1tuK�R�m�]�|���\�nor��p�L��Zȅ ͜#Ɍ�����2�����n�K�����y���F=Iit����->��]~�����*O��Ř��"m{����\K1 ��qD��{.(8�c�]�`�vҢK��&��og=@�(�k}����8k��7�����������.z����D�r�*���P,���Y�o�ɐ���Q�!�GK������fO`�`�
�0����)�&�3h�aA7��[�ަ0��~�K�^��>� �@lٵ!mv���jj6�9
���B�ü3ݹ�E��a��o]A��0UEw�~��p�X�7_vD`JT����(lW�� �F:�3xG�E� �~�n��ƀgpb��^%q�k_���Kǆ�K������v��W��'Wp�����J���������ڠ�V~�{�P��R`�*�bBq�f�Uⵠ\��'� OQS��|��aJ|k�@o2�E�p�X(����y�M?^�A��������R诈�v��2��s{�@�GL��$�~9IJH M����
!5D@#��)�2u�ʧv���,�,G6H��/.�K���� ���R�M���衿�����_�N9���5��j4�*k�1�6B�7��-X����s��$�1�c�X�Z�ԫ���Y��0�S�} �O4w��)B[���A��`2���Ո�:D�O�Mp-;!V�HH��,˗����o�c�NJʹaw�M��;yG�aC6N��14v����lU/�7(3%zBI0/��N�z��dA*�cq�����NՁ��ؽMɶXa���"��h�`t�f���u�,�Ũ�|�k�&jؠi'C��q��/a3�;�߇�ה��EA��Xt7�ޯ����w��٦*�p� �xZ�	��S0�V���Љ�V9ޱo젙7H瘮�5�k��N�.CEU����[�|u�*����$lКS\>t��o ��������}^�<^�Ɩ�Z����!CG���<ә2p[�Z#�T�����M�R����a�y���_�'TD��q7| ���>����MRV�{�A���Vr)���z�(���i�*����O���t(��1gC.�\�f���5
/�>ff�T1e�_���>� �)K���'� =����QSn�EQ?Y}����؁�9aA�����?�����Q�K�v�%�K�1��dD����A+�O�1���A�zM;��M3��I���Ő�[�ؗ���Z�hx��>�����F"4�^jf�Vv�g��eS uR�|jG~��M�bT��V[�Y��?��m�vEo��Xr{�#�����No�U{J7go���xd����.����Jbrad,9n$�|d�3���m"����_�����_G{�Q���ˤ�{�p��g9������BT���#��7ӎs*v�e#�Ð�y�կ1v�k�K�\�l|58b�<�&Uc�%��9��,��,�e/����W��$r���'$�\HQ&<z-�72�zR�z%��{�'mT��|�D�Y��Q��o�ue�	��z"\33�����}^f�yM���%�u�md��Q��$��Z�#��^`;���&�>W��~��(����	��g���(I%68c�y;������EU���=$,��Ԧd�����n|wz�8)ݐ��	^���))kй�1�X�e+}��L��l�+�hhI�7:E��`l^�� �S���>7�#iէ�y�iE��H�z�(����4YՅ�(��O�XV�z��|��S��3+0&2b��jwF�&ݙH�����\�u��������Bbr�_�����;�+�l<0�f�rLNA��Ϳ�)��� �e^�N���=�H��U���)�v��X�C�׻�#rs^�hNU��Ix�K�P�o����wXB�S�f��t��*i7NX�n.�����u��[��?UA��y�A��]�j��e&_a�[�� ����*�� ��ί(��?��(�].Mx�9@6�����+�PRH�� �y�be!�(�?&��٣��RMIK�"����Y���[���I��D�$��4"�70�"5]-N$#���:4����n��7�J3�K�=캺B��}��*b������y��z�a��5�ʉ���ՙ������`3�T��9d0�R{��Z7���ȕ�0\3�Eb�4�
�fI��f��tO�)���õ�$�>,z��U�#�F�W����O���]�hd�7�TKeⷿ�Y
J�
��𩤎�Ơ�Ø��o�z�#��LS�ȹ��6����A�`qI��v5����Q4�x|��`g"��������u��O52�}���#���'&�7�@��`����7=�)\R�t�"�) )� �	����Ij��*�k�OD��ClW�jXP�rܿ����o���&
��t#ܠ��O��g}%9��L5�?��f�<���M]�g~?��6��{�ꣷ�l���-Ϻ�zW��8��9�1�5���*t����@S;����MoC���ۃ?H��iw��@��qVt=sEr��#e��j��N�!����@۹�1����7�0�,'6\ym�qbn���@�}�]��t��[��60���u��B�>Ȧ�?��d>�c�e߅x0�~�D��A�.-��`��ţ���N��� ��]'��~Y2���E�*3��}��{�3�F�$L�j���*n�Iv }<T R.���� 	2�WA}�~F���o�ЗW�0�k�/g��+�����p�u��R�X�[��,m�@�K�q�ṶJ���6ᦽ�r�iFߓx�h�0G�5,+�=;>J��MqvfqBw��,U����s���?髯���g�����,��{�e�&\[�bK�k��w�{)GI�LP��n�o�ـ���"\z$g[ˈΦ����Ι�'~i���z��#��}v�(��yz	�7�))\��1����^s^)�N���3�+����Fn2I��8qz�(K����G�0僭<���Z�5<��%��}�o��7����8DN���]��k�{�\_�g+��|W���8Cb!��|�(թ΁6�TQ=@n�S0��<p�O<}�A�3�15��8�`�.:Jr�:m���F�~�nn=���MZ"�&i=X˜]�On���*�?�*)�w�0?}�����B,����a\�[-:�Pb
�6�)�_$sD�9�����A�f_��ӧ�6���X���M��^^~ix��	@�`l��IB�jh$c�_����UϙUs�48ي�*�$=���|]
R 1�����K���
:n��W�Q㵮��%���=oG��uO ,�(Y-�舟������$�>�Y�漋��u���$�+ܚ���c��Q���y���"�+g��ղ� t�(�ǐ�51{�D*P��Q;�������d��n���b�B�D_��ozӳ��^K�d�y�j���\3 ���~��69��E��w��@Zqi\X�UZNG۝��)����H�ю>)p���]�� Z�o�2���I�6�Hv��Ws�S`���\��x���6f�MI~�UX�$PnT[�b8q,��B���S��H/{r(�Ny���,���7&؏EY
H�������c
Pz�IQ��m�xm[W�2rco$"(Յ�T�32r���% w-����^