��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� rā�SZ )����C.��&0C]�-��[�3�-���+��պݣ�k�J�vo`�A�����f����u�X���v�=�а���]Q�Wۿ�߸�=_Q�X����j>��Zw�K��SvX��ƥ.���#�����Z�0���#7{��\S$��@1I�QX~TQ�E��db����۰� ���>0�%�9�j汈��}��1� ��2���h�G��SeY�a���	'<x�p��k�H`�H�j^y�0�s�78+���ֳ�`�R3dW��_��{p[�?$�s0��#�zS�_��bH
�c�p�IL7]� |����Q�� ��Rr���=��E즕2%�����`�^��l�q-�]�p��jf��Ӽ-f%H���ȳ�>��+���M�71��4_�) 3�46h�rb�J�W� k�h~K0�>P$�_n)���5�r�j��W�J&޴o��$>��6��ŀ�;A~<6P��K�~��f��*I
�Z��}`q���ApC��n���g���3��-�іrO�mF���,�$��@�BI�q�}��Ȥ֐����î�䂧��@������U���vU������ �T#K@f�㯁����|95<@���+�-�)�����K���FI�k���*@�m&���
���ma1[�2�u�I�\�U�yu���o�|��2����;�W�W�}P�K>%5�'�8���׫=����k��,�t�M�0�8]q3���N���GvZ�#z�HM���f5�����;�q��Pj����H�L�}��T7���z@�o	%�PFmy�lc�
)�8yIf�o���Z�"4��r���o�6˦��)��"�~���6��}�pY���]��
��K,�	���1D�̹�@��$���(_kk<| &���x,�u��Sm��Fģ	U��U9�k-��c�KU ��1$k�):h�����!�Έ>�l�B2A�V쉀�#� o�Aڐu�Q�%`��ܸ��cb.�����E��&�Ѯbz-V*�E���bnjۜb>W���z�<\UlA"���i��J��Xj݊���	p��k��1O:�$w%�C�\��H��U���Z�W��k�B�E��d��/���|�0�=o�g����/Z^����X@�N �Y*E�M��j��Ʒ�G��V��$��Qhw-J���,�B�����>�n�N9+���̍�)ТP��yw�~2�]�4�E�,��$&�_�������%�#P� M����PA��[�Z]�ϒ=!�ܠ��T�X�`2s��gq�D���&��%�?�Gy���4E��[4�͹��*�r�S�Q�����!P<�g����j�m2W|���i�:�?���_7��[�@k��v��I�������,��u�T�䷏Cë(��5<-�����8J���R�[{{l�Ijt�d�	0�:�K���}�� ��@W���D���&�b�kݿQ<
�d�dl�\aJ�n��En�V���pT���u!=��$�Z�
���Ѭ�!���w�*�����
���1���}3?Dl����i](6�~Y�'��z�h[�C�;���[�K*����z�vAU԰��Wi�q�->/#��'�e�!2���L�Y��GO��҉g�@��i(��rt��Q�OyҖܡ�:+x��n�+B;�U��i�Os�Ȝ�H�`��d��$��v�\��@�\�����
��N���K��l\�ϐs�)O�)���6/v)����DM	�h[�O8���,rpl�ۨ��������7n$Xs7޼��%�`Q~]������U�p��;�����>8|e:����q�Few�wյ����F`��]�h� !S���4fᰀOe�0��{�����?˧���h��#��|���-�$TЋ��G�i'5(��ښ�<d�㐜t.M���1�4�!��hi��ϊ�'��g�;�����+�ߎ�/Y�:�VR����ǐ�q��լ}��Ĉ������[����������/�F���gDhOtG=�tl-|h��s���r8Z����CNu�R!CM�7�*I߫
h�����º� �"�6w3A�1Øl'|D>ަ�(Vd���T�=�N�[W�Ů����.�Ȭ���O����ǄR�m���KA�J���;�1��|�s��0O�	�IHu(wH��uI�&�Ǡo�~7�	�2����+���P
����F�~�5�I�(��/J��s�1���\L~�cR%�@����Q�|H��
iʁ3-�z��rW��Ͽ���5�D��XM��>�Fd��Od�vP�nu"k��1k^���Ҙ[������K��ǟ�	����ѥ%�~`��6�`�4A��Gʉ���63����A�ML>%�6S#~�V$]�f�k�q�,FsN�IR �z�1��*+5���V���!�|��f����F��wAʀ4n���V���G��3,=���/�(˪�.s1�I�%�Y-5&�>�*X}��X�^ᔴ��Z�h�z!`D�S��1$p�@�N �_�ω��S�k��T�
�aW�k@� �:#4(�0�gkH�I*� O��}����N2�K<d=�ޔ'2�*��������]XDk���,�c��{�~%:\����}�5�Y�MlOJ~�ş�$���f���I���`h8���o���Ѻ�ϴ��F��)�δG���A���}U����2i>�'�2-�:�۾[P;'��y��Fx��/��"�^�]s�������X���6ٯ`&4�����A������8���H"~����������7�12-dt����zL�d����ŕd"��I���l��L�ύg��xFv���M��n��C��iod�=����w��`{�P��V�d�	_�X�~u9��#.�h���j������Sϧ�p���!��,���%']��dPѥqͣRm`W�藙vwd�R�ˍn�,C���=���E������hظ��R�CeپA.�]j�|�TԂ���m��T�.t�8�*�8��z8���Pi(dɱ/f[~<W�����ɂ��-ѿ�n�g�x+5�ws�R�z��B>,��D,46U%�y��*�[�d�"�4�l��\zi�MU���eE�R��Df����Jξ�pcv���O}Â����e�g�����eO��7|Z�cͺ۽�;~�Ј�o[�7�6�L��C�#� )�������|��p6v��+���i����u��ToT	2vU6{��q���o���o���\�Y2H��G�~�"�<��*�1J%��uȡ�1��{y6��[bˌ�h������	#pa=o��&os�
nPH���B�vz���/�� M�/�.n3��\g�m�}��r,�m�v��:�����l��#��J��ڨ3iJ�����0߈�~�Ra,1&&v�*�L�s�sO��Tёn	�LF}q4>|�as|�>�Va��"L��!8��R���k��/AXӋ�My��!�x��5�1�ȁ��VRe��w<��y���E��x���t� �(��K9�c<h��ז��_�!<��\�e2
ףh*zlXFB肹�y8���Y{��]|�������Z�vh����@J%Xfy~�λ�`��|�!L��Pu�G�c���(�DO�$@���<<�Ms#�Ln��|��bEh#�|+סo�:��'Z�:�f6Q'±PN�����*�-�#����@��1�8鋁Y�G�E����hk'�Ɨ�\FsN��1��Y7���Ee����k�Խ�7a�y��7�#�6�:�]@Z8�rg��p\��ه|��?6:�`����*O��w���Fe�� v�Q������jCZL����|�>$�*SQ�p�O��b
�}	�T���4����-��ل�x�
� @��vxdP	�5�)6��۟��w{���Ei�R(6��խ ��T��"��"�v#L'z���v�W��Ć1���J$��,VzV���0��8gc�;kQ!�D�Z����YjJ�Z�1:�i2�w��{ ���)5N�ٹNǕKjX$��-�]WKYa�ke���$ll����tU�k�@�^��un5Ƣ��@%�?'���4��a��#�'���j��c}UH��g?"��.t=�T8�t�y�		+��a��Z�L��ßWb�qK2�YC��^��p�U����v�p�����sս�8S����4�#i���-	o�a�$������vS��o.;��D�:���vE&��*���x����`��-TPM�hL��V/�ȀLC��t��cI�����,|���W+��L�˂�hy�CmKc�<`�8�vsk���N��ۍ��:X�/1�d-�/.R1!�g��P�~���4F�D��I!wqd�bs�a6F����謦}�MV<����Q�?i�X�x����qa���\�]�`�(:�5�;JE%����)J���X����l�q;a���1��X�v;��Qƾo�8�dT`�9�|�]���%��{|���<؂J<k�~���*mOl[g8٥����aH��TF��\�J�!h@a9н�v!�}�r�n�q�T�Y�զL��&Z]�X`�M� -OM�ң��X�S|�'��#���42�������6���a����u�-8�Nq;Z6=�A�����Zyt��G1^Qw�tQe|9���RQ�Ρ#`����o�G���-�[��ܔs��!<E!Kmq��m���k$�7������9ت&�P.s�����t��������� �bo�y���6��*H�@������P}��?w[�++7s�����uW��M:p����+�,}��������i4ñ���[�7� �8��x^'�k)*� 6h�-��8�����Uh�4b`~`�`������+�>��u�5��OZnj�|h_nbJ�bɦdh�Ћ��O+T�H���M����)�	����~�M\2j�XǍU��9#K����i��ҕ������wÁ2"�YOě�=V�aV,��lY�H���k�<�'vHX�k �8�^)­��������԰x������+kes��`��Xh�Y=���r���f�χ��DO�&����38�m��"z��� �8�&MypF}����5�	� ^�����W�Wk�"y*6m���ݕYdQ���Kz���6���*u�6����K�h2.�I���q��j܍Ձ��?J���[�4��˦6���F7���AT�[|�uծ�]��`K�Rl�{��Q:�F��1(;T�^]�f����7[@ jl9��gL�i�)�v\��������α_kU ꅯ�NOe=G���A�p�j �`��L88�5���{�O��s��P5d[��C���S�S��c��]��_Ru�a�|	��ɒ^���YI�n�C�^�fȽ�ѓa�u�Aȵ'�;��ۖF\b���b�<��1&�|_�E�kRDS"����+�%�Tr^�KՑc���[&if�s���*�Hk-��/nA��\�'�v~:��@]M���0�C�R]��pw"DL����]SC]h�h�,t��]D CՉ �/�Ѽ�y`���F�Z�<r����������1xNl ��(a�Ө=o������bU�������$䉀3�����E�����_Wթ������XS�/�~a��4V�����o���'������|/�)����~"9�Z�Ҙ����0rg�2���v��X#��H4�A5���W�t��y sA/#���l�ۘg���Z+��ձt�����f�&�?5v�>4B�┊�T$�x@>) 5�=��"2��^*��� ��<���
M���_�M�I%;�����3��J�8�:u���%7�9"�1�a�(.�ܲV��5�����ACŀ]��q4������x�|a!�֤4��a��!��g��4.e���X�hq�P�!�K�Xi��1}2����\h� "�fF�q6K�Zx��>�`��G�D�7\Y`qp����^�;�+~���,�n9WE�,�`�0��>�
�A�?�8���	U�d��
�Û��ܛ����.�y���e��=��A�����J��DK�� q���a[���A5%r�����b�o�}���;�B\Ǥk�'�6^�M�vrƢ��܀�Bب�i	���G)�d�Uӫ5I�^�^5XZ~(s)S�k��.wi����^�wl�] '�Dh_����҉f�)�[���|^698�S'Ç����9�U��N�%��T�W��sAX(|��Ǳ'0���tS��+c(�ᣧp4]E�V�:I�.�;_Ϥ*_��:����X�=��3b��/���i���k�&G~����u&���&��pZ*��w�Ri��V#O����^Kq��y�6h5��!Բ��d���R��K�4��P��J���<��遷n��L�u���^�7U���>� 7A�R�1��͜V|�$�A�Q�a���'�A+~�׍D�g�S��M	&���M��\!]���<�ј�.�ki�"k���X<2���X���2˯]?��V⟋���?��$�d��$�">�R����U.���b{\u�<Ȉ�gS}
S��s���1q��t�E�[�?D�$��=����c#i��7Z��Un�ֶ�V.pk���1��
1 �
����>d�k��f!�A��[L��ka
\,�Y����T��ɁHn���\��
	I������R�u�vE $�+��%+�����c���tq$D�Vl'�B$���*����׃݋=kxݪ�!����v�Gu-CJ�@�о0�|~AԹ��GB� ��4�j
VJ��U�rD��;İZC���sr}^[v�WB�`zqfd��3�p��S�.-(w��uFΙB�t�V5������5L8�F8�&:�s��?��\
���I��ў�����|'Ku#��|�Z�^�jA)��ul�G���К-Z���~H�	B����	�!�"v�v��:�ۢ����
�*Y
p�����~(�l��ǒMlI��CqsY���텪�d��0-lS���*>mR�cH��+��R��C߈W�,��Vt���ֶ=<+a��|&4���gkp�eJ.GX��0j�]AH��b���+�q��6��� 1� Y���#�s��Z���1�p����Z��b�;y7�g��\u&)�9�����M7��l�E ����dg	�#��0���r�Ӷv�b���l���\�0�ܹ��3R�e4�7%�]���7��,3x��މx��P¬}�uf�OA�8T߾���ۂ@�۵`]Mfy�3�eT�O"uen�M{���m�M#�������_�9z�d���E%
�@w{���U�g��0�N��\���֚��\T��6�e��y���i.�7f����悽b/��G#����/Ɵ�OMM=�6"̜����q��,0b@�u�;+�녅���Z�����/C v~^L����l�M���ɂ�U���K����JM7�cebJe�7yli�HÿH��J�]o���`��@���cYlp��Y�@���t��æ�Z8��kTu��r�Y�cX���-�m봃FpFm#gE�&3��'_v�ѕ�C}�ZϪ�l������X�B>XAd�WH�O�/�D�\E����b��MŁnt*XH�|�������Z����p��Ie�Լ�����Jx��~��z[�0��fH��^����rE�˘$����G�D=����ϒ򳾌b*����i�0�KpI���{�_����5�Y~a���&P~��]��1F�6Z2K$	���%���}��o/�B��I1v���<�΢�0�K���ʭEv��\Um6���g~]�|���9�|��0�5	L�?D�Q�KB\���w�T�T��Cl�p�GjKa�l¨���4f�7��p���o��@f�vvE�T�r��GQ��}�?^3��,����A���>TQ���+���.t}� �}&����:h׽
�[V��ו�o�R2��V�)/�+��ns�ɡo�꯻֖�]�~Y1���tȇ-PHX(�y�=�dʯ�Z0x1#6��*�%���h���(�]��w(\L,�� !6�}�uQ�v��{'��;�SZ�k�v^�*;��4�ò�~���u�B�dF� g�~��ke$X�Nv�������y��W���0�X���JByg�z���T��n|���j-Cx�'����9)�)6L>���E8�J>����IoT4�CJm���z�F�����r�(֟=q�ƢU�x�����ƻ1�m��y�oz� ���Q/���b~�|�j����a�xu��_�s���ժ��c�\�t�@��nk�Ɉ���i�9�"��sX�(op�v�W$�D�ihv�Ѕ�j����\��͓��b9Xv@��I6g���T�(2-�C�?��Ý*V�G�о���D둨Rp�l���I>��`C����<'�^
��<38�� rk��Vuڬj^�e��ܼ��>�ef+8w�xV�0|L!'p��#�߽k�=�e�^X��<#�U��=o��wc':�{��$���)0�k�y/��Y������K��<]r�RHJ�,�Oġ�Y�"�:�?� $L�"�LY�s2�	��hi��$Ω�,�X�ܱ%} ����;����Z$�G�*�@��}	T
KMȴ,�Ahl�#�糇s
��n�.ɖ�;A���=-F~樳���:��]dv&p4�+f����s4���|j�9! �q@�S��p��]�k��-l�LD��l�޿�bMv �¯ ����E,Iur���sH,7�ztpS�8�yG3�|'�� �`9YFٍ��o8����F�OU
���?}��3vmqkZ#V�"��֜��i(��eP�7EӘ^d��^�A��ؔ��_p�t0)&q]��n�Zy�Mu��:�	L������a��EqC����;���"�F�]��,���GRl@"MQ%lp|���梮&xl���fNa7��d��tؖZ<�[����]Q	�J0l'[j<�I2��Q(nz��L��X��f����P�=6g䦔��UkR�2�E�vc�C4�c�ǳwYVEL6
�E�z�ύ�]!9��a�fm�J	���z�����i�=�M鿞2r��)�'��^H�<�(J�+�K�7�e(x�����:^f�TGK*�@���O@V��\`�]�П���/ ,��]������̅g��|E�=�s�
�����L�3�V�hL{��|r;�|�Z*z@��.���:���F�櫉�8����3��Bc0���*�|f��U�/����Q��rbx�0`�z7��_P�e��Y��t�!	���is �u����@"v;T�rؓ/T���ֶr�Y'�M��m����,���6�e����7�֬u{���Rꪜ�gp���^ҝ�`M񢆃�"�㙁t`,���7���T���3%�,��nݕ�p�y��e�����x�B%����.(Sia���* �x��ƾ��R9X�B��:<�k�"Z��U�	`N�r���"�q)Px2��CbZ*�+B����������[w�$�� W���ژ���0���&��Q��y���8��o��k���o���8����P!0�<9ςk0�����f?,
�w�����*��"y�j�K���k�A6#�X�Q��^׺tz�q�1.�M��x%�oTI��|�|7l��صa�P���tOKH���ǁ���:�/�'i&#�A�k����_k<�m>#��yN].�u7Қ�8Uk��<��l��X��Pp�s���w5�^�z�:0r������C5�MK�Vm��!��t�6K]�;٤�ͧ:�k~�D.�J6�}���p ��A�Y�V�N���4�Y ���*l�Rĝ@I�?�|�M�
�ȏQ�iƖ�R���t
�?B��d��un�(
�����u�oIE��+���D����z-jHQ��]F�-���%�경{hb�bhZR�7y�Ѝ�%���{�;�������|),�Z�>g�� a�_�r���Q/"�'�Ģ.�XO���H�y"?[�C�j&)��$��_����o�Zn�bWqprz����;VS�O����/~�����5�v\��[mF���]�z�m�K�N�x@�f �ED��DA��Ƌ�Gn�ۮ�H�eog�A�0ڥ�g�<7��ÿ���Uc�uHY?F{
�s� �Y���x	>#u��5h�N̆M����'�� ��'H�<���8���6��d���r]�s����@,Ҹ��+�º;������C�� ��z)��~�ڣ<�r2�H��i%}"C+�F y�; ���_�W�Y� ��)*	B|a�t�h�`�����N����M���jZU�&I`��МS
y�9�p��G��:���מ�
b6�κk���ݛQ�i���I�82gƑ-uN�:��C�SRdhi՝x'Ku{$�Mѷ-�4p�g�Dǒֆ�1Q@&Ro���}��h��Ws��RT�2u1�U8��ҮiE�ڞ$�a�g��mҰ��Liɜ�U�잳S���(E�f;BctJ�KB츓�
���Jh��ckPUϝ�(~�6����$|�6�r.��k�v�+�Eb��73$3PO�3�Q(�d��h��E���C������D�f:�W�H��(jCg��:�1��S\�@n!�j4���c�JS�[����v�v���sg�_�L�D<��޲��&�!˿8e�i��hu�mq�~UyG�\���"��ð�Te6Bl�a8��W�Q炈�|��3�U�=h&~�,r4��huJ䔵��/�y/iSp��D�츑o�|�Y�>PW�c	j3�u����}>��^����q�.����Kp�w�+�RM�ސ�0g^���B���hK��j��F�~�U�ļ��@R:f,��:o#k�f����3��:X�]����C2�y�X����6�?��0@�l!$j���������iŋ�N�r*t�!���k>J��O��ྦ��D/N�~)��y�W�	а��g�+���KсV�8�ۡL��͵d�
�c��ES�H�k� d�9��ҳ�U�z�V�����WMW�L+.��K�\����vĳ��4�X^��˴��_I$#��V�uL�|M�A��-��F�d�Y�4��TV��}�_;��1�-*y�I�UU\�]�1�<�LǮ4K	9��45=���B��Yjf!�T���J���\N
x��7�6B�8���s�;��1���=C�:�S��/�j��}N#�U�2A���8�]��s�ԏ�:�+�,�jW#�{���>÷�;z�_-�,��Dk��y�Ĺ���w�'��pWh����3k�m��t�Ðhbg����5�E
��.�����,��/���Z��C��)oe���jA�V��y�o�1�A4:�0�3��+�j�cs����>�vć[����Olќ |����{sV}�s1F=��m��H�T":�{���İNe>�:o���2���E:;�ߍ�W��{�!GfE�	P	\��$�B�O[y����⼹��#ݎ�Kb_����0�ǄM������*ӭ
�F�]^��ѣdT�d�;����6��w�;�U���~.�"�$�gxaQ�ͣJ��͂�^[zl*��`�z��&g���������$�mP�Q�sH�/����*R6s	��p�I����|�q��%����^���"/։\�~}������Q^�
\x�F��x�#2k����_*l�ֈy�q�XD�T���Вf��b����y���0��F�_���+wц�,l��*�b^�M�(�����|��:B�/s�S����0�n�ܸd�!������I��/�$����`Zٓ�݄ohf���
��B��;G��ٜ�?a48�#<���L�n;`��Y;�^_�R��+䊇����&���X2wGe���ƥ���2�������(o�f�}Sb3�����Xg�M~j!307�>3o�d��3�6�*/���~����)�q�������ZN@Q��bΚ�	�7%^ѕCl��{h����M���xu��B�w^����xmj@���KD�4/���0�cgK�^C��_�r�VZ��U� ��l}eM�����ç2cI����.��aР!��D�)W��l��� �o,G��� ��=��XY����<���bNa�1g^��SC �n��J�*_>�?6��܅���%��J��B��g�F��j�t��>�3:��g��f��B�g�'[�)=9<��5�/��ş�@v��*�%[���'�W}���i��N�TE�����2Ƃ~n'�h�V�]yg�$���dvdm<i?f
�I���#x蕵q�������ي����'ʒ�)Utw��$��ӠK_�q��q� ��CLo�����.���p_���Wg�b3���"�,Gg'��@Bl�������6r�B<�8�?ন�#��[���jzS,�:��'k2eoJ�(M�c���(�x�,�p��g���+���cL��ǖzL�y��+�m��e�����3Z�@l�S[�f�׏177@����d�-)�rxL~t�0�B2��|��s��$8$W���v�K�����u�L�< ��T��T�!		=��Q� Q��V"���iT��9۟:��ٺj�ϰu��|i���l�5�=TJ�D�x��y���
�n".��j�K�>�`�����h�UF�h�h�'��ڝ ��Xi1+|��z�Ti#�י.���
 <������D�g7_azn%�7Y��R�*ڑ��-�-��ۼ¤��2��v_�X��/��$,@M��7�UG䓃+�nF-<.k�씙��Ԋ5$�Y<�s$��URu�����;Y?C��@D=n�q�(�1���nlO�Z�
��$�W�f�ho��;�g�{�֨��O���dEn�ؐ�y�φ�^��!�������0OΑW͝����D~�Y�$[ �_@�f��1B�ĥU�������,s�9��*v
��|>���O4��4C�>��33ɔt�B�N���%=����張�W��	=y��wKq�Uj^>>���YL�۞�ZW`�ټ����Dj�0O7�\ma���q��)Gf'��_�,����k2�+t����7�u�UL]�F3t��qogr�R��D�؜Oo��	f��C{<���P8�t�ٱ�	%�%#_d#[`
�����i`��_�&�\��5��K�,�T�O�5�Dx�X�Zb�U�'��2�	���w��#=1�=�Ô�G4�E���I��q��a�Y�k��n�"_��0J��8�����U=ǺČ2�@H~�6cY��	Ί��hT��n���xxP0h�����H�gb�.��"s]~`�Y�m�։�RW@��4���H�ς���2����"YM��kx�$�貅˹��7�e�F5����TQu�;��1}�3�?��HV�A=W��u5�g���m��nJ}�v�<^��2f�f�-.�QO��
l7��k��ӐZC�d��1@s�E1����Z��ZA�	���,���dqb���J������g�k�wC��C�m�77��OTȷ�U	�/��������{��=�����T��m�W�,!Z��ǵyL�ݠ�χ�=�� `�xI��{QD���+�9��xj�(���AQ�~�����DX>�"���ar�v����r���t�%�Vx=b�?��6��"���W��'$:�-mۯX�k%�&��fS�EY�|@>���O�F��L��Bn�u�J9$��y� 7d��8oF��w�F��YW��Խ��^}ڋ��Xz������ܑk�'��kuV�B[��y]c��3R�x�ɪ�j\0o��( z��˽��h�^osϯ?�D��������2}�Q�P��H�oK�����r:'�M�u�&<!�Ӭ��j,[��XG�5���-��9DD�xD��U���h��ר��S�q�`�fLU\��at*2�5���1BHq���,�o(f�d�#Zu�q��G�[L�e�掸�� @&�t A��X�Y}�h4��7�������`�P��^�"s�jW/5k1CD��-�t�'�1���ʡ�_��nՑ�Zc���$����!�ǅf8h�ziv�u�P�]_��8Z����Kj�R��a���	��Mݳ�|��r D�
(�1��q��V+��/ַ�������W͆iq��׻�q���i�0�G"��o��D|�/���� 	5P�iaz���b}@�t<fs�:F���Z���<�n_��S�4�%�6;	�Z=?Kd�Ig�I cUm9�b0��;uQ@ޯ��R��.�_	���Reԗ��ۗIr���|}���)��7�aS�{�>;��*�;js�:���	ြ�)�+��R�zHT��,�-G��3�U,��B��a��뽕M�0�z���[�k���	�ؠ!�4H��Z��i�^�g%z�ؾ��x$�j-)b`�4w�cZʽXG���*e��ae�����^E�N��q*[�\sad�C^��ޕW��f�i*��8؉�X�hbY�V�3�g��l�*9���L�A��e�ە�A0V΢83Y1�jWWr���x_���_,@�iO��X���V�AK���W���,/�t�_��7�r�$�����û�h��T�r`����3I��me�Q�i}�c��e�z�B����<�P3�n�_m�ٔN�*vN����x��
����R"v�E�BD/F(�+M-�n,������D�l�Z���;�O����%�R�� �4���#���mZ�Ei�gJS��Xj����غ�sm���rq�zuɄ�^24
hL��}����w��g�2��$l,�-A�+ⷄ��
G��7# �ݜ�?�� �iD�q�[�ù��<	�lx�;�퓸a��DRW=�f��G> L������^��V:�]���گ��p!�1��F>�tMW�ޡJҊ�������m�����~����W)l�>���||@�ԩ$	� ��x�1*'��� !(i�ܕ���Cɡ�|+�@��KI�'S�R��Y��9}�"i�b<o�Fc�r+���޿��j�A�fN�]4$����G"��/��T��g�R�i�iB�#�dKAy23���a�N3& �c�K�0;�.ޫB����$�U���L#�*L�����۞Ƃ9�4�@�� &Ļ��7�V�6�)��$���!I�[0H�ߢ�F/�8�q��SD���ׯw���%�7A��tW�-��|�Va�IXU�Ӣ��O4_�E�kw<S�ns]^I���k6Y�ܠ����ɎB2=��6 ��ͼ!>��S���a���!��^'�6@��n�) ���:n�l J���!�_�R���`��ړ����q:$$�hM3B�UINi���ZIĈA�Ofp�(���N��eC�
�]�"���zX��,����w���Ѭ���S�p�-{�s	Ax&!���X�8� :��K��7[��b�@¬.�b!��QI�oF5��,��"\��A�G=2^��:��}k��)%uw�1�p�X��br�J�/�BU`�lb������(��+`Ҍ���Rk{4p@���m�p�;P�u�n�#�+۞�0�q�Έ^rԵ�)�?\_P�e�Mǆ��\P�����ĸ�1�dw��Jy��@�38�t( �M�0�e/=���dW،���7���h������j�����{,!����M�|��$?���@�<����;���	�L ��@���O�X��#�p)��[��t�p��&�J����;s��d�<��
#�W4Q���[,W��0n��<Gs�J�3)��Q�]��xe�f�IF8�z2,w!7�8�~W�g��yu-M6o-�X@&'��Bq篤��-��M�YtW������c|Ѩ4�����F蝬�{�XN��!AJgQ���>��<�0�9�F��i��ŉ=�)D�;S7v����_A�s^�h�:����r����y�xt�Y�n������|d��َ�Ef��m�z%w�����Ow�'��&����g�L��C�	!�f$�X���AX�8�Y�߸Dg2	�B�w�Ф�F�3���+y�;q��e�,�:iV��m$�ʂ��_tt���+�N�U�`[nc�Gw����=`�/��~�j�y������)�m5����+JQl��W��
�#�����{���I<�N���5�0>[�n�v�j�)���C0My,���c�Ԕ���2�"��7�o��(���`e���D^�9-�,����[�,��e?�b�Y�_T�qg��FԚ�b�)o�ڼ-j�u�L�
��|�����g�?���|3���޳�f�/;U���ɣֺg4J���̵~39��'м�W1Y�BL*H�A�^F�3��/.ۼJФ�ةJg;���4"O�L�cR����MM����P��h��q̨nDP9Ɩ���Lj���Y(;�*��(_�U;�J�,����=�P��w��cmչ�(_è�a�O�`==���j���g�xA�?�	cرg:G=�B&��j� p=L4_ң�����BY���#d�VG�<c���sH�pt����9/��ɇ���i�T��1{�����B�Y�2��!��1��("�3<���D_~W��� �.��a��V�&���lF��O.)���Ͼ��W����'���CO�.�ۗe1�; [߈2l�,.u��(JF�����h�`�Է2i,dXwH�{Nj_�h���b�,lͥ�����$�T��z��h����oW!������֢���*�|�}��ݚ[#0�x'�f�/k|P�����DDD$/{�A�*��p��Ecr����4�a`f��?Z�u�5s�d�O�n��jn�A�ˎ�\ɟu�1&���ѡ�^5��f��a���meF$�S�;�)��9���~G������������L�|��X�L�G��>*e8ǂXAd1_Q�-���U�2����`���6��-�����]z2�ǘ���ߛ�-�7�����2"�u���ae���ƃ��:Zq�e? �c���jg|�6�N{0����8ܾ�n�0v�ev�)������.x'�6堙�yYde)0���&~�o9�Z7��]Ti�D}��/H��u�3{�3Y�����{#��:_�1C�T�� V!yh�Q��W�>�ͽ��T����y���jpػ2��Y���f�.E1m(V�N>j�Bg7�j��c�ځn4@�2a���Z"��h�k�E���%$�V��!��Ί��9�l�����ی�L�#A�5',�s�?m�������-2�g��R��hu�u��	�e�A?����z,O����1Rk��"y��)�x��j�q�,��8R�N�WO�)h�o�:Kvz��#�����\�ĹO���5������جU�?b]�i}��z����e-�1�H;0N�n�Q�O!�'�XƲ�<r��ʟ᧷��)e��X�B#�Or�g��.r��ǽ�H�X(4.U��}Z�	L�ej��%�)�@��6<�x���Mr�Fa�{��P}�[�xf23��P��⠚�CY��Z��|�<���r��We'|U@��#���	��O�1u�f�ڐ�ow\[��r=m&^c�gAht�|�Cx��`q!õ��(��;~�9a*��ɰ�`�v�dp�-!�[AX�o:�w�9+P�'+�Մ�<�jO���N�V�b�SMθ_"�G�c	��3�#�U��Z©vN��*塅8�i20	���M���lYH�)>_1�tIo�����3c0�B�RZ�t�k�����b1O��ar �,���%��sF?���V�mwc�I?`���L~����꓂y�U{�
q@յ�}��x���kIݖ�|�ր.�0	`/�s�T-L'	�u���I7�q�B��&*�&4�����mk.��}+A��D��������_�!�{y �|˙4eb�\���|dD�f�6�0c:-�#���r[]���7��eW>rw/��wѮ[ԆWH0K�Z������`
c�����+�؊�8���J����)��!?�nX�.E���rI�?ޗ��pT�Q���i7��mH����<2�xʜ�c��^ku}h�5A/��A|�C����z�F�y�ts��7���"{e'�Q�;%D!�W%|�(����v�� q�o~��+�z!mp����_����ꁼ{�ۻ����J�(N�,�#�͞��`�a�l�L��I���l��l��?�dA6�1�<�"�ʵR�J����E���u"���txd�SLcou��F)Z��j�+n�f�6��'^s�z��zs���*�=M;��J��}*vo+�S']%t�ү@%�[/�?����[�T*�`��0c]mw��B������υˇ�T�簜��q����m�;�N[	����_�q��`^���Fh�(��p��SL:]�4p��xnU��j8P����
r6�9�Nm�2�-���GB�ߥ�P۪Q����ع�/�:id��Ap%���b�w��!c�';�j�a��m+-��tYH�gK1��v}�>���C���^�˨���zR�sV���1��>
�u��պ-R
�(�"�^e��$�����v����+�.�F���Pͧ��)#�pD��=�Cb���Z��0�r��+��Q=���i���w��-�ͩRf�(\ž;D2�<�q��g�'XJgv�^�}���=V��(�@uZ�2��-��5@Ӧ�L(���S
�/�,6�"��V��ُ��* ܊4-�;P��-�.�!icw%<��%�p�[�9�/��:PQH��9Htz]���=�Ͼ.�6j��K�6Љͧ+h����A{��r��u���R�_��)��ro�KzO9���E��D(�밅8�[�@���ɡͯ��[�����~TL����������<~\���Z��),>��"��xD�Tr�/�Q��U"�Kp>L�~N������}�(���u|O/�Y2�����YJK�6�Av�8﮻�}L^})b�!������֤]Ǧ�6:��ǂ�z��I��8�z}�ô��(����vg>�E������m�O�uuO��a�0���n�|g��M��S�>ή��
�Dv-�׻uj�=���m"�;����hG��d�"\l
�9K�U�!%*���5�(z28�7K�ڝؘ��iɘ�m��}ظ3��Q>vpn�TZ�\�A\�8��r�Y"tL*�u��'���H.8|m>��{�
:kBae�Z�3��0�Ir�Y^���b`��!U%���x�l��"���"�7sÊrC�Ҧu�kc|�������3Hh���S�'%��D���'S���;���Aҵ�&>�����h�M�U����t���!UU�P=@�M �]lͅy0�8�����C�p��g�V��2�7<�ȍt�S쨩H�|�	vo}�G0w��uݬ.)�X3� JQ7v8bwx�|x����l�xy�J�?����ŀ]�/����mb�c��H�Oa��{a4�=��^%PyoZ���L0�7X�U�����,؊��#�Q
�`���(�����A�2�i���L�~6/���J���J�R0R��OD��y�S.��>j��#)��ZcZ䩄�g�2���%>�Ob�hx�B�ݚp>�W������m�ɸW����X̓�����I��˞c9+l�Rx[4�s�'������P�r�H���'��� �"�L��/�'f[�լ �tF�#D0d�z� �4x�,��j��s?���7���8A-��m����"���y��`��f(h�H�-�8ll�9Ц����b��W!�.55 f�-d�s��T��`��A�5Z�8����&�  �1��[�w��ze�zp�Ǒ�9��}���(��l�v֌��п��eꔸO�he����H�MG�nzb5b���wx�����:�n"x�nÊ�?T��b쥼�v�ޝ_�������;Ҁ	���" (1�wDhߠM�Ϻ�#7�aR��Z�~K�[�	�tJ����M����g	���j�Z��KP�S�<��oT���%#g��>��gp�OO�K�ff3f`J����ױ��Sj_|f=g��;�gJ1��.}��ɸ~���M��zy�u��	�)3i`��@�2fV���Do��}#wF��5�9�V�&)������[�5*�s���"�m��y@ `��a�ƍ�0��:u�wnBA��� ��b܄z�K��O8�̉�9EF[M|(�R�o��
�D�#�As�i�zp!�3O�5�ذ]�1^HXZ��-�<��������D�-��Y������l_��))}5�)�/�	V�c�iy�����8���5�GD��/1kv�����Q����&T6�1_����>���Y�@�it�5���eO�]t�d@����b��؞�P��+g�I9i�~e�l^u@�J�+��������߳�2[\�V)�j���2��K���<%͌fW�*r��0����}+���V�������r㰜�׍7Jy�B ���o�V/�G��ꊫ��`�m��Gt�?`���C�������q�-F^ �#Gڡ�듊��Egr'��ǯ�B��8�pQ�,'D�H~�݁\�*=�]�'���U7�0rȠ_��׹L�հVC��RJVd�O�Բ�$P��� ���Xl�	�G��!����0�W0-�v�<�y��>��vu�]��h;�Bx�|7�Z�Lt�X� ���%�S�����
��ʿ{�8�=X��,�Bi��w��ʹw�t��C��B��~�J��_��D2�ox�$��1VS���m���,ɩ4gr��)�~C2�d��܄������x���e���$b�}��ت�M���lٺr�����5�^s�G쭾�b���T�s�2D��H��e���. ��׉Ma9��(���M�8�@a��T�˚��]��]/:����b����R�'(�����l��?��?ąo�j�D�
.MR�F��q�L����Q�FYP�`�ӟ�����
$�8q���9����3"�`�?âF��c[�N�t�Ǆ=��L� 24�V���-�mR?�����ChS'#8Ng�v�ה+*���/�u�,�ܨ�W��G9*��[����gG���o�~P��Ťrݎ!�\kBl�*RHx�����f{;�Ak����Z���V���x���%3C�����o�9U#Si�����FE�揍��WwJ��"�K�d�(|w�*�eC���T��Tk����ø��)�iu���<���b�q�����Y��Ư�m\�����yz?r�?�G{�"�G��h{��V.(�Tך�GH"pPo�?
=9�1�s�R�_ӵ���5�e����:��rSZ�I��p�h��Y)����6��+��?)�� N�h��m��ʲ�m��k6c �g5N;�J�7ž�M���C�F�c�s�hp� 	�ӽvԆZ�r?�?�h��E�	,����ɢZ�|�6׃�o��jkJ6�sphr'G�jf� ��`ٗ���A�3��dN�p�Xۣ��_�T���Y�q�X�����Q',O�Hϳ����F@rL�8�%/��H�ޣ�´�&������t~֖�]�)wǄ�94�V�:)�:S��ODB��2B��.Ź���F��\K�S@~�v�"|��X{�����A�b�<�W��8�]GB��'������5x��hg.5pq��{
ֺ!4��s�V�f1��"�۝�O��4�~W���k����VyH�os\OG8-]zd"�o�[���Qᭆ�!>�]��y�ʩ��Գ�	r�@�8?��V� �d���������#�Y�P�zZ�?wZ��z�,A��$V1��)I�@�¥3������T�z�l��O�z:ep1`Lu:x�v��Ӓ� #P��H���4�B�y��9�s�5de�U���.+�2��q�������K��ժ��̟�E��Fd�G� ϳ�_z����Z�N�A���S�����:j�z'�[>U!�q�.M<�#D��!ۿ�e<?Z:S�����%zl?��
L��*A2���HH�oI�[�`=�C?b�1�q1���b92y�\�=��p�RDPˀ�?���O	��=I�W��"�+jc;����z=Y�ĵb`i�d[�	�P^ �^��"&8Xs���-]�gh�oS��c�*E,�>%�MHP�v")����W�	˞�w@����(Z49�cYϻ�nŶ��O��Q�;�#n�G�D�������B��I�d�o� ��{�eaXZm����񷄃m,�&E$*U���e��;V�t��db�<��S�01��=�G<�Y���V�(Ҏ� N	�j�ܖ��N�Wp��&{w�[����V,bN�����yd0��}��R�[\�����+��?x� 0X���b�M�vq	W�69)-̳��b���6?�f�-ٓ� 9<B �O�I��a���̀X�-��-nψ�;)kE��k#���H���5K�"��т�٪=b���eZ z/C��b>������s=�f��*bm�s iq�E^�}����8���y{�Ϭr|�U�C��mV���Q雉�[O�٪�D�#�)�%}}:��g�(V2�'�=Z՜��$�;&���m��
&��>􁎇M�Z� \�7|��,
j���R��ܦ����օC-���skE��{dO��sfѠ�y�TzČB�q!Xܑ��᷶��b	kd/������g!���q����\�YO�i�X�,��\U!v&���Pj�H������<�W��E'f.��x/�/�6����$H���Dzy)Y�^M�G��j�����Er�K᱌�4A��[$ԑ�?�3UL�v��F#{��׈q3��G �~�C�9�a��z~�����]u��"0���Tu=�c�6��R�DFH��I\�BL�s��X<
W���y��Ǌ�{�E��]�ǩ'2����dce6�&�:�&������RS&�M�̍��k�蘰[���~@�AC�v[#~��ß%<8y���g�����J[������&�YH�Q���]�ئףd�L����b�^�s�?`H� NV���'��F�)�5��-Hu�ū�`�6�(�wk^���<y� On=�Iʳ�/�U���l��U�5�U��@$x&
�O��]��{�l�ɺ�ڇfM�P�7��U�ͨ!P�����X*�4�B0V)c���4? �,�M�/��n��Z8g����<��j���ѵS�>sM�n��$�@���gG����V&іt`�����b�SH�u�	1 A&�/C��.�1��Qa�&�H�y�G�|l_|{�UYq/��X��*(��H�	C�����P\�#5����.¨��ϻ�Й���e����3vҧ��#��:�	Ý0��W��24֊F����Uq��.�@��kj��;������5#�,�pw�Ƶ�o�:�$Z�����p�o��߃6�/����
���33�@��r-����-9���Hl%��}����� �c�@����Gc�+$e�����E��L�B�Mj^���Da�.���T ��F#�FcQ��!�ٔ���3����q$_���8Z�Y{��@��[1��i��-(2�t!:a������[%�e@Ds��T��ೠ1.��DE ���N3�kZ:�t4�!~�H�-J�f��Q[e��Z����_�b��������+LM<�^U�[|�B�aD���D����ڤ�
_Ĩ����� O�}7�vjKc�w�K!�`fjc,�T��������PO%���͢���ɪ��������j�KkZ=��d��S�f�$���o`>D0�''\���r)'ї�%�;x��e]óNv��O:�k�mL�e#
��h4YB��x�C�O�Z���Y4Q�Q�����q�(���;� >S�Eu���ڲ��Z��R;'a���Py.��1/:�/~� U�at=�6��������@�Ћ7��O�c���:���;�I�~3���Z��ZG�D���QL3���s�|��<pʠ�s���d4�t�@��3<��tdZ� ��K�j�$�\��c��Q��JƊ�ZC�\ų�����������r��a<����;|ܛmH��H���Q$s�ǧ#u�a,��1;����k�l���r�H�P�<;�Ϝ~.v��[�8��Z|�f���$��?-
�T�8��H�{�'��IV͜��7p�kǫ?��lQi�a��u���"�;�	~z� �N�ȡ��k֊���L�[���"訝
�]�W4xWv���*)����ŏ�*9�2"�`�a ��KV9-��ޏ����7x6]�y���h���6�<7ca<9Tg����t����.9�u���da�i&m(j��XM��1��Q�����땃<�j��jщ�p8���
9�i��:���ܥApn6����m�� a���4���<@��mǌ�Xop�QEZ�W6eSD���h��T��m(��2��\�+L�Z�ZkF�K5�%D{X�����Dg��TQ���}������eNuQt5�K��t����D�Fr!�q#P�������)g��=-�0�Q'���2�Q\(�L ��i>��_�(Ҩ%�$��������a�}�*!y��k�U*#Z����@_�����eD�x��u�=n]ôXy�5�YR�mD5�t<��'X�E�RU��)hϳ�}���ܓ�������ɛ.�5�(�8?������a�Q�_ᚩ�M)d�"}y��f�T�E�R�>R���q��P���6����Ϡ�)�B�6N�G�i�����F���3�"xG_7��(m�>nn�D��8���&D��a��Ә����/zk����+¦����앩h�j��ѫӠa��UA�Epn���x�1�bfq0��e���<U�$`t-��{��(�?�c/Q>�Z�o����^LW�
�>	ǈ'���� 	G�l���(D����(2Z*:4�a�q����|�ɂ�<�n(�܆
G�O�ŪqEN�Ҵ�[��[�[8���lψ��)��QHd.�e/p
[K�|��zOB�N��D_KN�:�� ���z��s���Q����/����d��d��*��N�ٸ��.X�������\wD���:��ck�s�޷ư�ub�P��٪���,���.��I����^�}�_ ��fU����p�A"�� Ƿ��&�j,�!�J��L��NP����h�	�E�XH݉�T�ztr��R*���%(�;�_VZ��'�]q�dQ�5T�rњ&e.��]�xg���~�!�$�jy'�ϡm4��?�:��~�#�]U��ũ��{i�����ՖQj�#S���Y^����_��˶��$����x�Tg�
Ȣ�G��	����_>D?���j��U���X��g!WB(!��m$���#q��Cd��e���^��K�Z��$!a�ug�p�.����ܶٿo(j�eR����Λ��PU��2��O��IO�kh���=����9~���jG�%$���z�%���J��k�F��S|�e-����͙�07��N4'-v��n��������rA�,��-�T��J3ըR�������H\���^Eߧ��l���&���<R����nQ���n(�v���F�V�at�z�����%�ؿ�ûi��t��zR��U�'D�<���a҅�d���>g�B��?��/�]\>�R�������y!�:x�V������y�E��nx�A��4]*<��Rt�S�+c���՚+�J�ʜ���(l��*�0F+�'P(Tv��I�����v�j���I�`�Ou:�T�����	pZɑ�D�M{��)M����Z��r�N����O��E�h�x�o#�P�Rpz����WYNQLb��N�}�t��d� ��Ia0k� ]��_��+���8���Z�4���޳NG�H�"�рI(��8��P���d�$�"z�z��)lǏ%5L-Ȇ�q�+��`,�1���r%��ÿ\3�07������yE����{�S)a���TB�6hP�q�j�T�0�VKxDf)g�cm�� o���DʩF�Ip�}T���Y�6��[�4�oO��>B�ۨS��N5T�)jhQ��(58�s������]Hc����������.K!l�=��Cv�%�k1 ��8�&��ƀ0N�nJ6��A� vnj�&Wm��"\/���x����z���-Ȫ�_��mʝ�9pǠ�Q�H�M���r1	�r�
|�rl�Nu����t�GbL��D5�W��s��{�aq�s��;J1^d
� R�b"�2�ԟ��f�g���{�������z�ocҬ��)���|�ў��KmÆRR��J��g`0���4|֠o� �y�rD\��k�R[�Ww�P����~���M�.�PWJ��,��i��ߒ�Cn��Z�*,�!��*�N��r�5W�]�D�߈Ĺ4���/�Oo%�q�`�4���L(T��$e;����"����sKT�A*�,�&tm{������8���|G:R�$��̗'��%9ݏ͸[�
d���*�ȓ�%+���|5��u��J[(�Lk)�#z����n��x?���ޠ�ܸk���i"ȕ���u(HK�����H����i�(��%�������4ka�8�fc0`:�z%2cm�"����w����ڟ�\1c�u8�vÓs����}��}���J�f4W���'�d�}���Rۺ[k�[a#x�i1��H2i��p����TX�F'�� 5<�����6MX�&�U�������:V}p||�n$ԩqJ�O9�SWLq-��n����)?,���t����$=�X�پ|���:�ʊ.$���b�j��/���E@�W��(vV
�{���H
d&�~��6������8M1�A]d_��L�3~���Ϙ=�A`��̵�lcN!Rx�j����+��5�@J�^��CZ�;0R����Ȝ
��.p��p"sgzAWw�s�M۽^���.�O��X(�#�42l�;I�$��?RwB��ی�����<ͣ����_@�Ǿ=ס(��D+���C�zK^����b�Ͳ�2MӚW�������r4wVf�����.�[���rn�f�����!��{�U6�≣���=���~ �̠�^Y�&�l�������P<��	�OT��{Qn�����+��5�˶�t���
�a�Gl��04�١�"0��.��P�hYf����/F��o��D��"�,��.���q�$T��k�Ĝj�='�	:�@�0X��0���<����R&6Z_�1�KA_��_aS}��C��?Y�WqI�mgz�E�M�qdR|�C�O��G{�F�w��m�����J�~�����\Y,�jr�1�~L!��J�U�@+��o�`��|Iۻ�Uv
9(�w�
��#�ʇ$�����͝FE\��BLFBo��1r
��oP�/��ѓ�H���Â��K���6��c�>`b�������0dSM������nȂarג���FqW���#��[��)���~k�Q'}�ed�l��'�0M�X���]�/�/��'��*��QA��SSb�é�)��L�"3a�a�r�7	�5�,�u ��L�q�S�i��2��[�:�T jkjS�>�^<=�q7����Zݭ
i�{X�[=��Qc��m��������20�c�̇�A�! ,�����߿8�/��#��x�Wz��O�)�#g�d�[̙/*�?6���v~T�Г����{����`MP&ֳ�,�j�NV�8|��{�R�I���[�pd���KAo16[C�]&������\O�D�5�+�J���U�	���H<��	���O��R�婇}Y�{�y~��M�s�o�X��$��(�	��ǯ+r�"m������y�YҐI��Y/�8M(��('u1VA�c��0x܀Y<0�,�P$��)�-��NDwC�v�[�14�<������o�(u�of�A28}r�G�U�\�sW��u���@kusL_a���.�A��2%E���Ő��k$�L 5M��W�L%�:���QͭxC��5��`���s#�5�/&t��ȫ�H��s��1� :�.��	T�\�T�l���"|��U2m�خus#�Ѵ[���̃����)HS�I� ������~p!@S��q�L�E{�ʰ$�,!p��8���4�������0��z�{	(ً7 �#`��Ή?�����rL��LTG�X�=��
��|�y��CQP<i�#��jr��\�*�#�P#qB��0Lk���]��O]����:�ҕ��/N�����{�M��{�9��Y3�y1;�&ϲ&|�e��QHBF�.�W�����C�#y� ��4���#��~�`[[�>�>�ӱ��7�������H(��d���UQ
6��px�i��dkg�O6n�%F94x>��Tm���Q�*1��g0�v��[9������
�b��&	ݞ����Q����I-�K����%-Bt4|Q}�qJƚ?�{��o�_�f�x�M��ʒ����gZ��H�C��'=}Y.�p$P�i/Ϯ�ޝ(8=��N�e��u��BFN���K��+!D�-�q{B����`b_��V?�kԾ�t����<�k<�:�l�ߒ���
��Fk�i���h�"y�Yq�0�ޞ�aT�~���8��5Z�"z��y��ã�uCP,�_�Ӱ𩄲�>ؑd����Ԧ�m��9k��|�nX��`�(�1���̸h!m�%�j&g������m�������1����?���J$�ܷ�;���q0v:�j��t�7���F�h�,=&�	������}Cn�3����3psi0H]��U!]<`��x��_��>Ƣt
.�r� �_�˘���< +�gwm�k�7[�$nQ���iӢ5��B��L�
RRӽ��U�j����0���g����K؏��Q�z�]U�R��%!�vRG�O Fk�l#yȶ�Rퟀ֠�<c:Xd�0ߜ�J�1�i�3�������<�p��
e�.D�E���=�(�j��ͭ�V!؁��dǥ���H���<���"��v�=�����yu��Z�K�zc�:V�1 �K%(,l�SP÷�f��Z��I�a�`�TGRX�$�����8�+U:�i� ~�N��=��$k.+�R�x��R6�Ht��1b�I*�"xP�YTӷ7�>e1�%8��	�nB����T	��`J	Q}���vPu�`��HW�zH�*�q�%
��J�:�x��.��հ��GU��b�ZY�8�5�>���W�{߹��$��܄"q:���K+度�7�Ƈqڀ�� z��!ao�s�����k6��*��F .��HE�%؁s��4�ؾ�+��c�vz�?H��������_�� Y�j(Ϣb�g��ŷ5�GIS,ZV�O�[�ǧ�&�4&E&U��1Z˫24�d��CX�1�K-ff_������G�N��G���,H/�D�	�yc�i�x����3 o�5k��X�����t���^�.;�[��}� ��p��X ��5��#�Dl�ϥ\�0�����u�}�;&�@뺍���H�u���(�t�!qovxP��,b���a#⪼�M�,�2)W���6ȜA�nP4z�]X����*	ë�����=�@9Ua��P�t�"n�˜��I��oD:��+i�v04��1|�c�ʪ��)�	���F���`���VKԗ�%]��Gcn� $9�d���n3@�㹊��LF�	+�M�+z߯�ݐ���۽#{�,��>ZH��?~]�>M�\�塙�.�QiG��	^�ڬ~j��Do�S'*�b}�%c����N�i�=��7�	'�	k|�A�!n�����&Q�����OF��]p������<#�V���M�V�G��=����
ɩ�'1R�z&�zI�3��SS��LaA��*w0���>��4�Nd]]$딬�����R_@^"��b�E�ֺ)���|�M��o>c�J?����O�C𥉉��reJ==�HP�.���&�0 �W;{�2�����YN�a�ګ��Y	��SVX�p�f�����T���'% ��/}�[XP�z�b��{G!�*:�}~�]M7���]�[��F�e:c�3.�IM��n�|�,��pV���2l�B �Ƙ&--�����~�`��qV���@;<R�0�r����YOM¨ 
��
Wa'0�
`���%�����K?�-�B�#�I�C��ȇ;A�UD�g�����Sp�!]C�ʆ�pn��}��<�:=Ǔ^�� F.#��0��Ȩ����ti�W㓷�p����Ю�^�k�%�Bc)N5;�z��/��������2	��<뉫R2f�/cf`�`͞j���_;��^D��wM��Z��'�]|�����W\=m�[���|i0���8�"dl�oa5��is��q���=h($(Ϝ��J�x+��&��!c*e ��'��8*Tt�+��;�j����ǐᩲ�M�ϋ�����o���0�� [tG�λ���}��U�Hü��xQy�@�5U�x�����y�@x��x�����-SU���_Z�ѝ�7���[-h�j�!+�H�jR:'?=���<F�����Q3"d��0�]q����VK�2w@?��A��忆2���W���O��^�6�����b���llQ�c�C��i�%^�)���A�&�����b$���,�t<3�3�T&Hq�\حKV��b��S�~Z�	��$S�t@����X�,Y��h�/cV������T�mç4�2��0�m�t~���b<�;]U=FNz�zb�e�KߗQE�W�l�,N�g�V�Z�K,��6G�E���v�L��h�?��p=Q[�T(Z{'f���뭇�H2�dT�x�ԫ���=�a�ï���M8jbC[�����K	#�W�9+���;�ۼ^P9:R�I����?A�ǧeǼ�7,��s��'WQ�������ƈZ��ET�)�4|Q9�z�w��rc�eb�ӥn�h�L�=����&,�4���-�_���
W��l+!9���:�ѝI_�&�a
�m3��{6���m�E��i��w��N�9��0<a%�y�Db�"����K�������f��|��o���L��wV��"�G�'SzAt�|%�1��$�����y��ʼ]�|�� |�����=e˼���r<��s���ef�}����!bE��&9c ��1N�iخ@�jՍ�-��mup��n��8�� H� ��O����/�a�/��-|<#Z`�D�j���"���t����B:�����}5�#az����fQ6B��3���+���1��dpt����gYs���N�5#ɐ�J����p7�?����H^�M�Q���k���qa�W�x�ѵ�������r[g��o_ԝȟfS"�Ԩ���׫rʟvUNr��ѱ�l_����	/�;�_rN�ӳ.�������s�"��R!N��D9Kb��ͭIM�S���+���>JvR����K�=a$�̼�����Fq�ם[p�\���}��ge�w��h?�<�$g�7߯иJ�\���I��Y;"yK��WT^yKp��=K0�	]f@�ڬ�nٹR p�̬��h��0���U+B���ݝ�N�?�������T��L�,�A)�������ɠ���5�}�?��!�i�#X�Whk�)�X�+}$��n�?��rMi���9���H�������.������~��&��k'��O��z�Oad�ge_Sg
?v�|T�Cr�2+��)2\��η$�Ѿw)�NoWIS�jv��>E=�r����~�"/�j������Z�+�D��.��E|8�.�����/��0t����9��SN��e_0zUQgj麰N
�Q`�(��Ǚzy� W��F��C�[��x����H��}L���t���E`�o��iO�]D��Ǐ�RO���c	4�ݶ�筚�ϯ>\��-@�)k����m�1���֔M:Ś�rG#K��f�A�A�ܙ��V1r��F/�ֵ����:���3�m����L�jW�u�7��'Ӵט�=>�C{�J�@U�qʷ�p=$xm�eG;��Y���7��O�.;��+�qϤ
��rb[9�9�?x��\͖�1�W�i2����s���i��p��?3g���	F�����r�ibG�"uk�&{�N�#���g�.���������|�+$��^�L�����v~a2Z��9�AJ�;�|S�XI�PsCz�什iE2x�s?b�tDߘ0���(��*�2ÖJ�r�lLZ�扡[p�����+^���i�3�ZZ�i"�D��u �����l��c����/���zL��"�W'�6A������I����y�7��<<��_Y�$�2v6��7P�+8���u��nh�1�84W4�'���[�<���Ւhy�q��z�W���ܣ��[�ۊ�d{Xx�oW� B�Hav!�0N�5�������Вw���a#W'���~���λ�����3�%�R{���ca&Rm�=��a�������e3R���������a's��[�
���؇h�7w~.W�te��,��V�i�f�F����
��h�s���?'�񈧿uJ�w��J&�g`��#RI7��6�0��:IG:����=�����a!���y�4�1R��Ӊ-�mS{$�J+�0
�������p����`䦺c��a��Ay�n'z�;���_����mH�ĳT�����g"��h��ps��W5�d�2�b���DRm�MLm������V�y�OB�ZW�4,��!~���L� 2r:�t���+��6ݭsp�$l��䆌��.������%���H������]�ɪRrw�Mr�y�����_�����7#���Q�q��;��=qf���F��ճ農����r|�<b濔�JK��(��v��P�����;-�$
8:j5ԉ�M0�������o�7�!pJqg$G-+����z�oE��� ���ߕD���qW
���	
3�~�1���*�cL#X��+�+��)���ph�*;�ϥ���З$Y_�"�F������I��]���K_�����^ߥĈZ�F오���iM��e���/��[��c���rxyKꄴ�SV�P_�ä�إ����zUn�MQqrD��jh��צ%��IтC0v�5e�.�Q�6�(�Fe)�/��)/������ͻ�Hy�@����~�Ė-|�x�l��0�n6��2��`+ɡTSH&�J�&��q ���D�X�����Q�{ppσ�7p��E$DÌ�Փ�x$}���P��TM�u��:o�o������=���vc��,FbTbI�βũ���w�bJ��G�%�q�o��O��{�sy���L*�#��)@UU�`iN炇��͆x��YN��5��!Z�룰�� J��J&��9�	4�k�'��qe�|���H}�F�Ů��V�pC[��RL~>v�wV�}TZ�["����:!��P��E=�Z)�>�R����_���d����jG�L"|�a���8ވǚ�&��`wI��+B�ŅeP�]/>�:�-+ƕ�+�y-���B�S�-��+�?ߡw����S��O{�}hHW~z��Kha���s�)�2�?	<#gQt�Jˆ[�<�ñ:�	��,�	�+B|���H^L]	�����]��� Ө�'G#�Mkf�x����Q4��u���`"�*i�FYUPG����g���������8�@�DF�C�	r����G8���b�r�����1zԩ�q6��Wⅹ�e�3�]j(�b�A^l#�)��K!�D$����G&�G����P�7��@^����m�Ltu'[��B���)��Y!cҼ�bOXS|��l��_l��F��G��W��~5��!O�#&;IY�ٜ�^%c�,�#/Ӳ���ӏ��ɼul�%7��S���ݍ3��'�"��D�-��<��e�a��T%����	����[�{�˘4S��Q��4�k���k�NssyJ<���E 2���ʒ?��v���w�S#R���ü\H�r�NA�|�垞W˾��&�/����mjs�j��g ������>���γ�Y!>I׵�{9Bk7BE]�Vj��}���Y$&�!a��~�>�=0�H@s�{l)�x�l���PG�_�F�<�|��!e>�k�-�!�&=��[��H�@�J�K�*���p�C�:�M6��