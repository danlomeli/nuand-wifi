��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$��7�4��L+Q���+2�"H�������v�ao4��	�u��=��d=�>�iV�f��l0�Zs��7���~rM��U�`���e����K%�u��ݒ-� rā�SZ )����C.��&0C]�-��[�3�-���+��պݣ�k�J�vo`�A�����f����u�X���v�=�а���]Q�Wۿ�߸�=_Q�X����j>��Zw�K��SvX��ƥ.���#�����Z�0���#7{��\S$��@1I�QX~TQ�E��db����۰� ���>0�%�9�j汈��}��1� ��2���h�G��SeY�a���	'<x�p��k�H`�H�j^y�0�s�78+���ֳ�`�R3dW��_��{p[�?$�s0��#�zS�_��bH
�c�p�IL7]� |����Q�� ��Rr���=��E즕2%�����`�^��l�q-�]�p��jf��Ӽ-f%H���ȳ�>��+���M�71��4_�) 3�46h�rb�J�W� k�h~K0�>P$�_n)���5�r�j��W�J&޴o��$>��6��ŀ�;A~<6P��K�~��f��*I
�Z��}`q���ApC��n���g���3��-�іrO�mF���,�$��@�BI�q�}��Ȥ֐����î�䂧��@������U���vU������ �T#K@f�㯁����|95<@���+�-�)�����K���FI�k���*@�m&���
���ma1[�2�u�I�\�U�yu���o�|��2����;�W�W�}P�K>%5�'�8���׫=����k��,�t�M�0�8]q3���N���GvZ�i�+ C�e
��Ќ�S�v<%���q��e_��
�k�夞��>ZO7E~��5k�TW Aod��eE���G���ɑ-'���?�G$����ќ����8ɸ+ 5ʗ���l�d��,�J�
�^�3b,�����J����#n�zK����z�&��;|�\�^���'e�W�����">�w*	FO�Δ��v�.�3y�0L�o4X_��T�A�{�n�aDv�(��@�s�:�
��^�؆6�2���8����Md����p��K=���(d9����>)�4(v�]�T'��( o]O�Ct�?=�]�)6J�;AZnKB��b4�C������f��;H�l'�5���٤�&��GA�8�;��Ӯ�t�|��I�3Y�OF�68����Z�9�R+{��!m�9��Oկn㊼h{�@��`��iX |5%&��|0�n�
B9X�`d~�"o-Y����2�Z%4b������T�~�٢Aʣ0����B(� ��ˡ�"�s�2��2���2H&	F��L���p�8�x�*�L��c�&ل�F����(��[{�=���BS�ϑG[&E<�]�J��{L���OS�2m��_�*���%?�Nr�D!�2}�R��?IK'@�Q;�
�ʽ��9]H���wC�)bcx�� q=��M#,w4�Rw��4����oWM�P��Ӧc�>�ތW�^טm�zb��qf]#�� 9��'i����2�q��&���MC礴g�>��k����i}���9��Qj�o@�(ܕ򃒞����Y�*!����,���d��%�q�a��,* �;����W��&�-E�mOx�/�o���S�+���9[�\�=�����TM6?���К<x��5FU@"z��K�
J1.o��7�=��_2s���,��.�=ӯ������=���O>��$jO�w���>�p9S�|��e�Qn���̘x0y�(%-_}��9���%5`�������n�U����H�*9��Dv[�4�Ͽ["^�7��u�_V�(��8%�L;���Y8�H�a|�c��/�z�_(� �R��w�dy�5�45�[�C��33�������CS<u] ��=���hf��M(�g"b׬�t�E`6p�z��J�pC�ԥ�m=Z�QT�Z��W��
bWG�b_�cݯ<���C'���TbߡP�\5�[�f_m>����B����;l|�b��?�j�K��df�����4���Q�4�ї�1b�Y�$�F�q���1�2	�~k^C�h5�1��������ilDf5:�D/<՟����f�ߧ�
������I%�3�&D9o�k��cF��\>�!��2��ɹ\���ח��v!>'��C�v �>C�b|�W���,��/���r����4˙xH�l�1����HqmXi;CiLt��*@>��ו%B���I5��,I����m�����u��i�	jı�f�3K�2m}��+j!/�h���w���K�ۯ�4Ir\Jgzm��1��l��w�N��S���<z��"��훏=��{��e]�Xdd:�3�2��rv�A���DU��{��5�f��B�a�P�zo-��}-K�Xn�:e�[�9����A}ltY�t��O[S�"�=�P1{�h����a�'�{͢E�O�n79�ws7,�8qE�[>M��0�EUf�&�P��9�k�a{�1DD�`��xY��syy'�-3�g��b �A[TsF���Jn(�^�A��u���'>$|^m�F�wX�?����݌:��~I�m6*��~��D?����g��pKU��>Z	�+����@� P]P1�S�ﷸ�0�����a@������&�Ne'<�sڳ��L���p5�7:�y� ]��f�szs��=��\G��sU8@E�t:���/ʆ�&�oU~�uS�s�7�nB��ػ�����L7x���V�ҏՈ{�qEY9��q	*���65�^H#������YI(���K��ò:�ܙc����q$�k����9&�p�S�R���h�6�a�i~x��Xuz8����+� !5��,.rT�
1��Z�v�Tst`�x�t�u0?�	�1�vrO����VL=���o������qz�E�&����HWb�܌�_�e��,��)��+xRs�� B]�ʂd�i���x��=��ʶB�8D}�v���a�$�*	bS���s8`�]���Pl���_Vf)0.�uQCm�����
�W#_���y;��Z�f �6�#�䘍���\xL�}�3�`"1V��`������,?#"v���D��+^<��&�qJ��	��2�F����U���MC545�+����;�:�Q$ =��*�q8it��2D�9�t-�ku�#l!�ʰa�jJٮp��[ ��	��|�g$J����u2Y/:��n��Қ���.e�kM4�G��p�p���?à��w53�j��}Ur���yf�����b�C::�̈́+��	���a���N8���%��J^0��ܵ'/�{�rCE��InZ�3�=&	'�>��zf��6y��T���]_��C({��2A���MK��:�C�up�1ݲ±�T�_�( hLjT����/h~���o�=���0�:����O�r*9q�q'��ʺ՝���1c`�)DO��eX��$f6�o����Kp�b��|��U����)6%�5Rd.F��F�{�u�f��Y/��������{\.�S��P�$���H۱ �wF�����r�ʕy�벥���/���|9�M6�VG�$8���X���>ԋ-a��:ov������+�o)���j��������\���
[��,�@���fM|�ծFW�&e��� ٤�<��y�t`��Z���sҌ��&vAJ��<i���|u�"���T�1�"}P��	�햸P|�Gc$��x��.�9��	X�؇���0�����ʡv�92H�?D9PM�`8�C'Q�-aU2I�ҩ��7�389~۫9X��%)6�!�|�Ǝ�!찁�� +C�F�XShtU`IG�'
e�76����5�+����c�h�M��A-�����3�H�!�"���+";�o󸕓0��H3rR"��Xxyd�z�N꾸����Y]Y�����1�J�p�H��޽������]��d��'��OXApt��VvJ����l(�\&��������V����-��ǶB*��Ne�
l�)  u�O�;�_��,�0��f�����$���s�.l�������`6p��hy[���L�_?��N�$�����)os���J��ͧP'�w�E�����v���s�km����1T�l��o5��8DB`���=Ҵ���}S���2��),��T�=s���Q-��m�K@ذ�T��P���@�&qxY�D"f�T[{*<9<g��Ő��~�x�������e����Y8C���H�;+�=��Ҽ�� ϛ?_2m/�wc&.Ƙ���E� G�E��5a� VA����݁���]m�Qm{�E%��m���0�QQX�D�<	���[$����i�wz������S�Qͤ
H�K 0�.I��y4C�*��4�#��n���ʞ�H���ڮ�0�>����^P��ׇ�d�~_uG!�s�,�4n�k�8@��.���0$bF��5H�S��*I�!���,UX{��pΐ���@�x;YYX�%���R����D��r�&͗���7����7�z��"�O�1Zv3��M#P�_��_y�ozt�"�)t^I��Ο�J��4��hJ��� !(1"@�Gp�X�
"%TE=�G�Pw�u%��S���;�vkw�x���R��BU���*���|�F�y9��:�YM�&Ǿ���	���O�ҳ�w�v��t�V�`���B�<�x�iD��x�/7�6:��׳ɇ��%҂��m]s.x�������`��$%X����rȟU��?��ٚ�}�o��g����"����)ќ�/���m� �~3��~�sAN��l�Qv]�~b3�m��{ ���4<�-Q��q�pR9�Qy�K�y2n��D��g�u�]r��;��|�5�v�}�\��{���q���F:�7�M˼�PkG������ы4;i']�H����~rl��h�w�cGX�;<�Ӌ�Kz!ێ�d�\�"��;o:P��U2���)(�U�y������ ��z[��B�,8/��2ƙ4�z�i`o��ߙw�6�\N�1���#3��Y�N���O��a��[�s-�
u0r�J珊��%;c�~9��~G��~�)��UmFS�v��d�%A�(LO�q=�гG�����Z1��$0�T��L5�6o��#��+��zs���y��Q+7���}$�0:����F$x��|��}|@����?ü@E���%l0C��NJ���"���� H!\����jF�.Tك���`s�Y֙�d���)�ӧĀ�_Erm��ε��-e��Ks!(�d��ca�P�5nɦ�h{�Bٳ�t�R.�����5�0;��2U�����D�o�"9[��9����:�t��b��
�؁�T}hV`$#z�W���6ٖ�yU��ԃ���-���#�� ��z�=� ��ڧR(�tVꠠ�c���E]B�������C���q�L͹kd�y�CL^��,��ɜ��4>@[+�h�7R4owkOrx�OU�F՜4����F��}I�s2��P�b�Ɖ��^2��42D���,��n!�*�KIA�$l���٬����lcA>kgi���X�Ά ��b���(!���d��NI!
�]��,�"�����tZ�MN2��E^u��r���SCj�&�'������Or�dα+�����;���o�/�:s�!h���Y��6?��A^Ɖ��_w6Ҹ�@��G��	���+�����lz�d]Y�h-;�F$K�wSO+V\N�����P���b�8�d�,��J[<FZ�����k#0��_xJ��`f���+WQ;�G�&9`�%��;�)��a�U>�o��*��c�do�=:�=���H�=��<�R~�2o�M;;��d����B��n��Ag��ܐxY��$�� u��S�w䣿��=-s笋O~ �:?��;���Lwg�2����L>��m�W���ຸ+��y�E�ʅͽb=X"�RŲ"�ׯ=��1���X���-"�I�q��5K>؄����N�vN)�*�q.+c��80ؘ��&g�����L52ę-?�bƱA8��6�_�;㉲P�Y���ä��xX������@�q6̲�0����'��g����!�*��Jd��Q@����^�\���$d
Q�
����B���l�g(˵�{��ж%9%v�.^Y]FE�[M�P�u�ژvj��o*��l_��|1M�go�/��Ξ�M�2�~J~h���J�/�r��͠"o�
���T���?pv`2Q�9G&��Z�X�*œ!��̒�̧L��x�β4�iU��N��߻�&E_���[����ո�/(~l�ذ`J4۬p�>���߸�i�iƀ�3���%e��i_����6�"ǖ*T��1�n��g$�;!*\�j����s�\��D�d�OHp��������v.��*GZ�)��|�᷉Ǹ�bT/m;S��ܲ>��?�XeʕP�J��@PĞ����Ѱ��R��+7�F�}
8���!�־W��"o�� Nr�d��X�D5�x��s0�t�)�k����8vZ�t��&w�R�06{eگ�qd�&�ą@V���ԒQ˵T2s���Ex���!e��sQ�]�H��-s��=!#�=�c[��\p 0��4,jQ�tO��^�����y���|vK��n �<�wViy�ʡ�e,n��-�GC��I1E��e�Uq��n��pm%��O��?W�Pֳn�������� �݌�\�4u3�$������ܤW����c���N���M�'���P*��dtz�W
j�5ћacJ��¹U/�Oۭ(B��f�bƾ�N��[Ľ��A%�!?R�~|����w⤀Q�%(�*i��k��(�L�s ?!r�sQ��Ŷ�T�������D4�1'�~���~m��q���f{an�f/)J�
JQ|�,�vQ��L�&!��9|�5�w�g�zx	�c~0��N �1�嶦s��J*�
�K��:�O��^��]��Z���.�z~_]"���|��>����/�yLm=����c��b� ��f�l�@��N���XL�Y�4�<��=�;�^�"�㨩�%vD.��1��N��D�Ө�����U]@D7�4j�1w�?��;h����@C� F���~��>�hG7� ��1r���zZ�	d<M3�XA��������X2�-�
cW.���\�i�� �UDu �7�d�v�vOl�CAٖ��� �)�=r˻WN~�MH����w���¹��ji�;A������ (���!�.N�eF�6į�"������|9J��)�K_��ؙ֕2!H<��=̓����ܦ#��/w�aCо�]�v�ܱ�	}GǙ�w���f�wE�ܚ�gǛ���q��y�&y���Oڦ}����
Xfq�@׻�Y�_?�׉�	���n�Q�|��i<��"#
� 7���wڂ.��Lu���7p�ZP����HK�g�Zh�� ���F�)�<�D�"}2\�Ћ�:9���w"�ݝ��l�? qTU�ԱN�QM3�X����=Y�$��T��x��V��9���^P��n�^�� C-n�w~2�7�=z�r�Dzqn
UKhS��a'�?�A����Ӎ�dU�\%�Կe�1����w�C�3�����e�kH�SM)r��&G��$�����FH�Z��7�48\ш��.�<`���x�� ��T��~?5s4��o��v����V��
�:�����0AK�{���-X-�!h�����mڝ���{��?Z��k"%B��!�7�Ü5�ˀgX��r2�b'�L����s�˖��ͷy�z?!$�٧y�~526'SPh^J�p�M!=��CX�ʛU���(��0�[7�
�����6ٿ�|���"�����2��{p�ƪE����E�U�9�1d��:�j>��f"'��)sK�\rV��Ej�:z,BZ�:�S��#�Gl(������$T*����&~��?�N�'�
@3�K����)F�}�#F�[��w�/�t'9y{CR bK�=|}O��o�ҧ�B��hNd�EC�0@��z��jf,9��L*�%�}ӵX�7LO2/��VW\ۼ3q�Q/?A��D����J��:��m����-Z��&�b��E0���:�qס�l]W-��{S�S���%�(�?�SX
�z�y%s9�>"N��m �O�oy�����5��|p��(����p4dq��p��U��aM-���"��dЅ�4���������r�#I6���I|w�¹sR����Fm�WB+g���^�xԑ������\4��?�p�	Hm�����QjOҨ�������!	Kc12�Tm���3�ԁ}?�pFۃΏ�V�`O��Nk+�x0"�W��U� ������*(���u����6�q|��5�\�չg^��i�����;�e`�h���	���%�촿��"V��a')w`��O�����K�)�=��r#�W��ϿYϭ�fj6+8ƶޔ���P��#�c��-�;/�z\X��[�}(��+x.�TT��":ӕ�Ȗ����,y�i5�>���@�-�gG<�t���4�Kh_~��7�h��.�Y�KnD�a��(�76sÓ�*���`*R��fP#�
6z����F򠨊Fg�y* '��W�h�W'���%- U�Ftp�ALE�R�JG�.��3Teb�� �W�5� ��8.���wZ��¤u�Sy�d��B���&VK����~WJ$�;�����������ņ�L���&��}}c]���x�h%�{57�;�`�{>��;yd���+�����Wg�(Ȃ�gȔ ��S�9�VD�O!�DIR%5�l�5����&�|ء�c�.p5κ�^�A���R�E7�P|��#��X��(
����CZSJt�$c\��`H���Ry����5m�6��~��lL���E������4�q�hX�B���>b׮վ4�5^���9��(�~� ���/���S��⪯yk�L	/����"��Ӂ%!%��J�]��(���~�Y�.����O��)�?TT��O��(��e_�? 2����5Ŀ��q���h��3�3�z[�K0��
m�`�+��mH��i1��>�aA�Rk��N��������$a��g�S9e���'J`��l�Z��#�O��5�$��"��~�1^��H��6�A�{κbX}��8&�8�Ї��0�y
���'A'�pa�ްy�ݮ̋�����[������ �^�4 ��`���i��x]�R������g�DB^+׾	�:� W���?��q�nkL����k�\���H-���n6wP�/\��ڭ,�"�Se�J����ژ����
8�đ��R�M��7��B��	�	���+�	@�j%G�ǥr��;R̤ؒ�ޅ�=Jq�Ԝ��a,R|J��*��&�;�bݲ@o�Nũ2�%�]� �[{<ح�c�G��n\��XI�M������	����W��,q,�oZN%��=~������R�Xm��F�K�``���/�#��1��9:V��G�|��+��ʞ�f�p(V\���Cተ�0x;��%+б*o����
$�������Xi�W��F�n���^��w�x,
V�8�h��֤�+-���R���giq��ڇn�$=������5>S�Ś&5q���w�IP���D�;N#TJx�v��kB�Y�q\P��D����=�'=q	��hƬ��rE���s���3�,93�����p^y?��=&�wA�����r���S��-�v��� ��#2J�2���*_����B^˭�$���3���+7jD����
��vN�qaiU�E$�^�N�{�r]�؋3��E9|�VD���.�9܌*Wƕ.]{y��b����0�/��e��~afa�%�t]e�r��B�Ar6��|~Cr�F �鱴sD��()�9�k��/Ȅ�W��qE
b,S��Yl��O�]VU��t�x{O���$GP$��tR�1<
�וW]�@u`P�٠J�T\!|]��J2=�/�G7�ǧ%����� �l=��m�!A�kKު˽�k[�m
b-Q�)c%�w���Ye!�/1ٿ������ag�����]8cO#�@%r�<ԥ�2�I3iͰ��)y��pUq����~;sjn���|��^�1����K���ai'�O�e:[Ö����B�DU�@O03 R�o�,%�H���$��{I�jl��!2��<`�5m�C�2����hZ0��rrB�����Q����ïm)�<CC-U����sG:���Y�W����P2��*�i���[�y�k�.����u�i�W�k�d�q�Lxn+/��ᨰ,�)M�OYPOx�p���/����i�X�Y$b74�N4F�����φ[�Y8�t�н�5���A�n�&��ND��}���Sv�9tz�� n�^��.�A��Dc���L[�n+˖'K��b�_���C+��d�0��������i��5�� ,��}�J48F�FQD4b<#��P�ǃ_�����O5P�j�>x�'ŉ� K=���oN�`eZ*�ջ���Yvg�!I}wS2�bgU��M�W����a��K@�^NG��S����G=B�����OO�Ҹ�8X�P/l!�2�ik ����~�wL��D����uƼ�?k�!��וg߶A��H�_#���E4�z�Ê^Q��D ����3���;�Z�TQ!e�i��'"7�5��M�v<?���B�fR��~]=�y\���Ni!E����B5p���)�c��KҘd��7���?1�4�h���B�F�����a�%�d}e�+�^�����sv@?�݆y0���,z�����(��(�LC�bŮ�kK�b��9�j�@��xL�}d!Pe@ſԦ�7�t������Z6~+I�B�[?"�T��k��:�Dbڏ'�ʷ9��K+�p��j[v�Tr�[w˗		������MѠ�]�$�!~@��ع�3�`_w+̢�Y|�����!��Ȑ��|��%���+v��S|��X�[8���@r~��%��7[�b����>)>���H荐�����A2W�Z�� v���5�%m��.�.�
$�J�{QE'f��s���TI�w\u&��)~a�T@���kNfŖ�p� ��f�AP�vyӲ�8�{y���T�h�9��W��闐�����_�\�u���xR]�@4	�ĳ:Bs�@�Xa���~&Wc���EE�d������3�����5vq�,��{Cq�}g�^�8@OI�=U^⥖e�OVA}��@_�"��
hΑ����&�<R�U��APC�by�H��dE��V��b�
~�BG�T�ļ���c�LRS���e���־�~����q�Ne� �D���pK��%�����M.�r���)ςΊےy3h�D��
+-Q#۪�2�b�"@Q���	�n�$4��ЙW�+`lυ��P�
����lH	@i�q�f��J�����tS�cM��a�G/c�Mځ�ZZ��6̤c��4.$�ju�� ��3�1'��:� A�=����WR�1f�/qaY���Qwk���m��l�ۿ)j����>��Y�p���'.�gW�X��GAYX`M�Inl�5�s�E���.��o��"7�;w����7$�z�p���$�����/�u�S.�*�,dT#u{ը�(��_q���}\h���Q�F���VTΣ�*�R?'y(����n�*~&Ug?�4���!�����3vn�F�R�
IQ��7����#ӱ�Ɂ�F.��ۮݍ!.}=�Z�9�	f~��%��4&�1�W���CPL��iB���sV2��B���h�4�^L�0�}��am�߬R�F��6L��LLz�B��wdJ;Hh�t
��e�<_�V䮃�j�}���<��:�k*dμ�<��⁁	�0���Nt5C��w59�h6oF�x�_��9�Φ"��\�*	�;<���g�T��N�y�y��bA���3R��Z�a	�蕧�5Ln�5P�\��$�UZBFkV�]v8���@��!/u�����'J�\�9Yz���%ޟuŴ=/}B�(`�<N����H��IC����(�H�8��r_3�#�e�
�&8HMu:�u���סd�"ܞ�~����\��'X���g�S)���Ot��GF[և1r�
Ш�&-"�\�2�l�..ǓpA52�4k�e���W�>gH���srcv���t���Q�䞏/�:v�,�����1��e8;����>	��X���9>z���lc� ��ÂL1!�4�wH&�X���$�h^~/��%2./ػ�QTID� yX�g�j���?�Pu{w�a\9���}v�f���wI��j�h�y�o�r�|]�İT������`0�P'UP���=�
z�C�\(����g4�ϡ�����\���{eJ��ؖQ/�i�u��=�.y�O��6��e`�mZ�V�x�B�K=�̋]�.�,�8�B�N�j�#,�;�.�Y�G��i�<6��ER��V�3e��+�6��U����XG><E�t\�ŗ���k�m�'���/��Ms�p���������kjn�/��	����e�#�iˊ;�<�e0f��sS�Cs�:k3i���=��6�-��'8���M��)y�b�Lj�9 ��ki��� ���9W�(;�S�A�v�(��`г����a/��Mv��D�1N{raD����{͊���%��#�M�K�ّq�".��	?>x$� ��3�u�ii]q��1�J��6`0o�˄([|�f�f���ݟ����:�\H�q�F��W�[���m����5r��<��8�Hm]�G(�"����k6�~�0f������-2��/����d�`�]N"��p�[r2�����L�@��Q���AZH�p�3i �pX��l�6�k���� ��"�E7��;�.���u��ؕ��Fx{��]i��A���h�Jl�%\��a ���w]�Ե��<�����
�^�q~2O��J�TK���tߚ�9�8j��	Nh�E��;�ס[��L��0=���s[K�Frd�X$�ݺ�7��[)�F_�Xi�S؃\|������[ ���_���~�d�(y��2|�yt�کi�;�n$ͷ[+qt9X^pn|l+��R�m�츂ĳ���e�D�Q8XS}��9���\X�|�,xl��S$��ɸc��c^��*Jt?��R�oٞAL�I��7/ZnfG����-�G�Q�K_����Vw�0A��#�]T�viV�!��}E���UQH��rDP��� � ���Q� �=������Y���s̝,|\�Y]7F�%���J��(���iu�v��4(��+.Ak^u�*SF{j���k��[}P`���n��>I��ecykc��a����k|��Ӹ2z��,�h�Z3�0��/B�/#��#6��t���۩!���a���$��c�F���K���"=��vu�Y��F�M7���.n,�n&e~�G�v�@]��p��Qo:ƫlVH6��ȝĭl/�|'��x��)�%��UÇ%����^4=�G)e�6�Ev֡Ē��ݣwG��j�
}��n����j��a�o�A�`~U��y�P�}?oJ`v�gP�]=0�<� Cz�"9���3����%�Z�2�� �9�"�T:��=4�ʱR�y������y�����gC�t6���
����W��q���]�o�EiV�y�eL��k�]��O2Dj9 �6�9 n�PU�3�r~���k�w�x��7�{���^jǅ`�_����@��J�N(C�9�1�C�ZX\^�W[
0*��\���y�2��E5j�m����l�@a�&cQ=@��o/�l�}Y���tSF�֕��V=��+�ɖ/�OZ瀿?-t
W�˹���`�A���U*$�q
|���!����$��H�]nE�e�8�&-އT��S	W$�F�sk&���=P��FY���$Ɔ;�V$�z]����᳙��&P_79m�#�+u�l���l�q��hH�' ^q�G�>-<��p����-�
�ݾP�Kԯ��Z:N�Ta�
#DC����ܭK�wX�0�T��G%��$)QS��!�A`B"���7����׽-ڷHRM�,	랎�1���(9840���έ�q�$���C�7�;�UV��1�eh�a����,�R0�ֽNˤ�\W���`u!���1Ȯ��l�h�lq���0<��x����Fq<�l�N�ȿ�ݫ���!Y�!�������:�2���sA�V�h��<G�d�w;�X��i!�md;�![J4�O�,�ܝ�l#��cY~]��7���f�1���܉$q�N�dY�:��ڹi�B`�f`���I��`��|~*�h�
�9je���.��1�Ӏ��(�X�{~S��^m]� ���*�h�P9r��G�R�/C�"�OM�[ڷVjʁ����O�$��Œ_c$�C�La�D�yH�1�o$C��|�z�Ӈ�A55��)�,Rޗ0�w߇�)�t}���e�b�k?!mL���T`���-�KN�Ig��j?��*�l��eP����wV+����w�Kte��(�����)W;���^�������6U�58��kB���� ܌��2� ��D���@�/����&rFo@�,(��.o>���5݆����
!��`����-��c�*BJ1I.,�n��}��O���Mh��/I/�L��C�$b&}�,`��ٞ�Wt��lVx{�l���T*�;L�P��K7�7D5]k}*��~��?�S|?�s|s�A<�d��	S���ο~q^��/r>`52���"��C�����$�7����p3A	ی�Y�p�O6\�ȱ|��e���!#PM�Q��B֏OoɌ�4�$Q�ݡct�b�����a^d\Y��B�p��}�_$1:��L��������<?��bw�N1�����d��%��"�C����n_�뒬q{��Lt�/-�(�2�oz&U8ۓ$G��>�@��H��_�LW18���$X(m�W����#s�/��4j��e���Ŭ�$]N=��R�j�n8���Ϭ��������	�D�Ҡ�Ԯ���X5������%յEm+�(��Bf�CEQ�5IL��2�!5=��:l<�h��Ŋ�*���4p��;�x!��pA\("0��qx:�S�T�{X��~�2�<".�m�v%�	��"nj�~Y������/A�̡޻����c�������(+���f�+M��Z5
z�}I �ir�� b��|���!%�Ȁq�jտO߭�ɄaD�N����st����9�o{Xc��{j��_������P6�G�)�ܞ��L2T�>�H���&�}L�\ �胃;��J��D	Q�g�|K�y �Rsq�GO����릖EG�m�pr2O�q�p���~^�g���W�����P��<a��	F�"�F���6܇�:�x˛'to�y� 
�e4��_�[$��0S�Ц�O�۔�3G�D^�^%󞹏���-��р>5�ãDʦ9����樤		)�"��i�2ګXk^�A/��Ѡq�Y���Q�N&H�i�.d�=�^�{�S�5?!�P$�Q�C�QYKP����&�@��Z��I��d���|�Pb9�c�Y72��d���Z�����d��9���a4�ud1���x7:��h�x�l�˳9�K,V�2�����ܚ�BSA��湈���h��j-�+
�ٙL<V{�_4�O�}�nC�r)kl����[���{��T;�w`K�]+�/�|j[ȰF�Pi�k�O�݈m�6R�Us��]�]�_,MI�8"��-�1�Ƒ�	�+19�u8ݐ�	�Vi��_y���G��7��i��G�_�APm]�Hԑ���[e���y� ,;�B��|���(�;"�6�g	-4L7��������ߒr������@�(�#���Cz���B}+�P��9�ME�}���vR=/_u!������0�6*��Ά�"j���w_.<�]�y%o�fS�N���5��-=��A��팠��ċ��2)�* �A!nq9T>m(���	+Z(��GtE�(jE�M���O��'��rk$;�)���{p����C�>L���50�>�<�6��:B�O2#M�-�5�� +ܛ�pu�\�ɝ8��U��(<|8(!4�ς&��0�����l$�r	Zc�0�I�x��5+�p� �PMp؟d*�Y���֨����ƊIk��PK��1�	�n1UG�[Re�{�-��g��ܷ:W����ZZRҺ>hf� �y�kZt����0$���S���&��t�uU���$2�
f�a����I+��F��3�Tm�q*�xu��~�sv0"��t.�`�2K�t��>�u�� ���P�U�8Ԁ�-%;Þ݂�elE�~WW	|�2j���׷��_+Ep�+
X�^v�<l4jW�h�r��TDWʺRAt"�"�A�v�H��i�*���7(V�����H�#	sQ?V��lO��#0�o*f>���{��;���V%��*I]VU"�aN`vl&g֣˲ڰ֌͸���8̫ۘ?w2q|���̍<n?9�t�(���k�
��v�<�@�?�fi�a�.$���o��)>�<��'���^T������	�Q���
�W�XU����κJ4���!u��a���z�qv��nd�Db��u��!��z=�@�a�p|��X�z�2�_��L��p��4T�a#Ȋ�����'=wo���),�e�ɕ�y%�#�PU�B8�� ���S&�j�y���"���� ���ʳ�W4�9!\\Rι�E���J�q9���$#n�á�N� ~Գ,L�3�/����D�57ǋz!��f����1Y���#t��?H)�Jj�V���&{W����q������� � G���3V�� r�����s�	��W\"��_E��C鋝��b'�&-/��b�H�E��<��ﻹT (0q�ZH柶1�_%�-�i�J\������j$>�I�E�Y�u3'�0 ��7��� "aZȧ��e�C)�" T&��aҘ*ՈC�/� �����>��Vz�~�"�&�s�mQժu(G�c�G�gvM� ����Vl�QM��@ߴ��}���D%-,3�X�ｩu����,��Jw�Q�&O�3��<c�6T�� D�pVf����9=�"�����Α���pI �p�?c�A{���ט�FF��e����0m��w���ʯG�高B��M��d��gQ4�{����&�fsy�3�}�7���Q��ƕ�Rw@Ǜp��q��`�� @���_�<��k\n�zZR�~�;F��ƻ�q!�g��#g�_��<�U뫌񢍝�竢�����Oh�"0i�ñA�q��ۊ�A�Ȫ}��~�p]�a7�ۻ�m��!3kLp��V�+�f������n�q9��0�j�����v����g��1�	����K�)d���E�s�H�M��tڗ�sݵŚ��j� nq�KqS(�"Mf�~N'4�8�M^�g�3�s�'惌D��Wv�!5��j�F=0%-�/��D��crM���!Fc� b��x�nS�W� ��:\A�A��|KR��-e\�v�+x�(]o��k�7��n�[���J�s��UG� ��kmjM;��`�1�$Q�>��g��z6���2A��]�C�|��Hz�Ң/P���jP9�K�u�_��B<�="�Jĵ�>3.��1)~v��0�_s�������(	܉#eK��!2f���4:B�BYa� ����1裝�,�q��(����d�!W���F�ÊqЕo�5��T/W{
�,�sc�����FV�ʄ�'�P� �FW6�����$̔��c#���<>�`��[�&�!��fw�L�����|�`��"kM,���_E`l����&��ad5�`e����;h�#gŤ�Tm~Ҵ�"lSt[9�����`���eU]jt�-T�#�#��|-ú\9H.F�?O\��������iW:�h�E�F�+й�S���|Y�P�,�x����ݐ/T�R����0���G�\�v��V���B<> 7�C>]�*����Hq�%'X�t4MV�Eq[�a��,�# #�����'�dı��mG��-R �����P�I��\�+���GͬR���+�B~.&�Z�W �J"���%�����І��{qx1���q����鮮��eLRc���^�܍��q8[A�\�ja/�r��ϑtvq��kE��2n�3�%N-��Ǯn�P�B�۴p����p`PL���C��L��T�#ӉE1$Y�:���z����R���.9;�4 ��ᵀ��V{�d�ۑ�4
ĥ�c�qB-��
9f�;[2/ڇY�Q�s�@�wݾ��ቘ�%�У�@����*h��A�iH]�)5d�����-�Se�l��u���K�
rR�U��Gj�EW��{�"�7l+��F7�x|j�)�\�z!4鳒���`M��ʍ��?}$J����58��B�Q5��G�VR��3����҉q��S��R�n9|x�gX6N��+޽�R��X�0c��G�z�b�x
��'�ˌZ���gw4�}o��!��	�/���.zWzv��?�H#	L�^�բM�����ή�lN�#�S~M���+����-��9�d���d�	�d*>��A Wh����gͤ1��������p4g/o	\��Fz�i���젢Ө�*>3���t@
�P4:_�[L\��Wx%��շ&��כ��.Q�+�m
��&����r�'@�]���� ��U[���VF��w4�oQ������ˮ��(��X�!�ls��p �Mv�>��!g���ǐ�"K�1I�;�O��TwJ��*��dHo���O6 �6���q���	 lU}^�u ����9$o-�)��:���S��KC�(|�<J_S`UFE�|�`��q_�G�����墵E��VzZW<�	���Z��R�u��|%��1�k� �ԟ�Ee�e�����?SFo�{��l`��K�ֆ�<��x�'�`��΀]Ib�C��|+��g3��:q���ˍ~1�����kWq��P��6��r;O8��ւ�c�3�ln'nn��	7���F!���p�NZt �A��ЊO(�0�D��n�MF����>�o�l]ݹ��׫ХǨ����sծ��<8"���)B��@� Z��s��3��� �S�MZ�Z[�!��1e�͢����z:��x�7�g	'�p_��8���S��n[I���؎��EV��_�A-�.)���-�w�<=���;�ၑw��R�ƻ|ʇ�<�Dm? v��'�1�t��ew��tտ�<Y�N�2�{�7��z��ͷc~�F�|f�Æ��>��ۘ��L#O�+�qMǕ"yU|��	~	R�N�	��P��j\�T �oC|6vA�Vwǖ�
�#,	�3�m�I`����%^+��)�{i��	î������nn|e����i�Ht���`���$�E� �r����h�����|���Q ��i/e' r�����3=���G��Ylp!'�p��.�OGb��	�{��n�]��#��2��%Ĥ~���f���Ͽ����<�W%j�@���
��C�j�w�7�����^Sp��d���3]��Ps�G��S�}&S�Ɛ����ٗ��bQ�����=�X<��L�X&���9�{׹�Xb�LR����]w+a&\���]g�o�}1x��1����_���M �V�E�����-㇌qG�����F����ˍLP�3�jh������N���D���{�S��c��w�T9�C�Z�U��@������H�.`˨ƑsK�!�s�ɼ�spl3s=�8�N����=7����~�L/�x�̅�'����ԅ����p�㚗�� k1+�㫘��á�U�@W��l�����
�n�����-j}Se$�]x�+$�B���X6�7Ȓ?����X3�<cu�]�ۜ!]�b�]ݩ,ל��`�����'��8N��u���bL�1X|-FC`}��bu2�S�DD�Pի���5t|Ә�ƆU�7�R"Z����2��n:{#����Ptk)�~C]?g�Ȃ*5�� B���rvxk�!<�2Y)� ����*̒+P��5k���ȫ��B�?��ND���e��U��ZݑW�ݝ��)<}˂º��48
�MNQ9IDe�� ΆUO`��Ü+Kl�������(����NǡGR{_	�57��9 ����3>90֪�,��Ń(
��- �w=GF����V��� g�Riy�Y(�+�u.,@&�0]b�����8w�@i�L��!�=�5�>�-��es���dy]M(��TvAEQ\�Ė�]���DXOm����ZX��E���/���h�X��,"��d�![	=��Z!�UR�	��5a�ado�����&�6�-^_y�g���&�	.%���uܒ[�Y�i(O�wVI�;��%YÄ��*�R�[F�3�BU��/����M��~���8��w�oQ�K9Rs&��6��]�@쉽���_��e#�j�HR����2b��L��Jgc���1+����*
i��\�@��p�_\)޿��J�ǃ2Z� �s��"�=)Գ�z'yk���ŉ�3ӗ�^ܒK�6���O@�i�bj����S�ߜz�_����>�f7K��i�A�o�*���&�����M�"C~�CCgwH��Z��1>�V�2u��W�{;�L�H�V���"�����\`A��9��.��S؁�������+b���r��#V`ʪ�{d�\�����,�0d��	�0F-����ĭ&�9��9}.�A�D�K���0�K����S�\\���E{U����M.��׏����,�0�w�t3`�7���; ��q�L�j��Kٝ��J&��c@���|�e*KP�ԩμA9��f�x��} ����~#���K���N��.����tB�����g��Rs�Q�i� i�#�\�h��ý��h��B�ȃ���O#��l��`ʆb`Liŀ4o��v�����$��G�7���f��@��N��s�A��Ht?o�$+/8c�Xp$>���(�
��Wi=�`,d;�����Ȟ�7�2�.��2�R_X4g"9�d%�3�kQ
w+���(G���E$�Yf�q�S){��m����օ��������W�>X_��u�Զx/F�UR�x)rH.{Bp��d����[����5��W���G�aEPݤ�����3a��qN¼��"vN
�v��{��^����_x|&3��FåLw�
�*�~�T&|Eya����9�&Ґ���i��H����d��t�t���M��DtO��QS�u�n-�Y�4SC2�Hk.�? �����ְ5o��fV�D|b�:�4H]�N�z�|�!�q��چSt���5 ł����E+��WC&�����)v#0CU-�;ibܹ��������$C�F
_��Zg�������A�o�,�KH�^���=6�[��MOq6��ϽV8w��B!����|��.r ���U��8�_���1V��~�۫���HWv@]��5���WF6���S��
��g4k'=����Ӡ��H�!�g�db���b����:�Ν{6*�Τ7��m�M��vnU��J�莃Z��`��uEӊ�H�75�vkM��
��3{b��^QA��R�!.$%�h��,���&��Bx.�p��,u�BI63H
 �y-K���]�A0�(����沛�%��zhW�X�>��[��ѹ�Vt|(:?�̰��$2{?��g�%s��)J���$����Dh�0��c� VU��BO�~�a����Y��A"G��%�_�X��Im$���`J���燽�C+�9%�B&q���K�&"s����^'R��F�Ԓb�iP�[��o���@\���\��v��sXMS���i�Nꮫ�L�l?����[��4ޘ?ȼ��G�v  �| G�Ju����F"ٮ�,#��q�߫����t�n�rr-��F��M!6��*��1�/�d�ƹ��O���y�'`�vn[`�&�H������5��.����y�`ҿ��>�dƔ�1��ٕ&��gA���bۧ�l�e�S�{b��4�l�K�c��H)�����K]η����5ЛPmm`�'�\_ٳB�?�V��l5��u�C�7wVV(�d@�2iTi��4�F���
�+�d��{��L?έ���C�ڷ(�gd�{����˴���Ɔ9`Q�$��5�t*���qX��p�t���	��Tm ��}W�?a:i9�������|쨚F�IR� P�^�����GA'$j����!�Ջ@tv�^�<O���(!���yx�@3��ԏ���@-�B��,��5�鎈�9����ﾼ�<��M�Z�ϩ4���:��ۄEۥ1VR^KК��a�I�r~�e�6�;>}��t�j�}��V
��_��??E*�-e��e�-)��ȷF�ق��(S_�u���0l��|��p ��Y�S��ཉ�3DX�L[WEqk<j���=��߹�|KA�-C�� ��V�E*9�H��)VI&���I��ߙH�ձN8�<��7ToR���l���ꭝ��<��b�I�������W���6�P�גw� 7/mpt��n�S��X�ދ�`y��r�6'%.6�x'�<��Y����d>�����V�c����>�Y	��w�qi��@����c�<�w���`�í>�'-�o@]����,�R��������3r����#�V�5�d�X��u���D����#��sk���܈�X7H{ZTqޱ����5�?���l�!��n���:�+�\��T�U�k�C������6!%�ı���vK(aޢ���-�P�54�bE�.
�x��y���>������NN���}��4U~ㇸ�#잳H�GB"Y+o��cB�\
�������H%��Dж޶��.���'{t��i�S����~��8D �6�gm��Z�� ?�ݒo{�(Y��hEǾ��������"U���*�Z}��GA|��`���d��RtQ�%��t,�+b�A�f&��I�>�}�}�	c9���5��i�;��f��b5�uR�s�,f�i���>�=���J#��$`�4��G>�&��}�8�-�xw�J�����7�N�:�CG�����MHz�M���ܭ���v����4�lhcQ��ʊ9C�W���m=6ť�Y;"hɯ?k.g�FP�֭Q�� p;��qh�i��M[�ś{������wK���_bn�ɜ��&�����K����.��{2-+������v׏>�ނ�u�I��^k����{�¤����^��>Xe�}v��L�Y�X>a$z�j����
��ۈ~9��#9�Ҩ�7�t�^�B��ʺ���!�^/�`�_�jb!�e8g ��ר�M������a�QM��P�����8%7�Y�� v���
ؚ����i��D;�5�A������W{�'O�ɇ�њ���WX���G�9�D��o�P<8loii�!<����҉���|��y�;�ܨ�e�Y�I��p��[�ي��_�E�:AvN��� �Q1��2��h" ���q�0�]^��溧`�i��Ƴ;zd�Άh(�\�Ȉi���ҽ�Y���
Ȕ�|����Q���@���9G�����ƈ�\8�J��]j�W�Eq��?e] ��BBrIAu�������̉) 8�Xj��Y���38ڍ��
�����X)�+H9 8��L�šY�\��g�K�1W�Q9�y�+��a��P^4̭�;���q`����>t8��ҡ����	8V� 5�_+����d�!{����Q�O��Q���b�A���{��l]k0륂�����eC�mF�9�|<A���݅y�8�-�>Wz��c�7�4���$��P7?��۩�I�r��pV�7UQ9�ف���o0`����̯�w��In�=
�i1�G��R�~V�"t���a}l\�� �}{
��Ć���>�dy]�ט���L�߇L'R����q�<k�h��F�r���9��_�p{�\&I��,�+��V-�vwq���.���յ	�	�&�al8Dc�i�3����`�3�bQIRU��3uZ���\N�:���)!A:��.�R��qϐ�3�j�x��\�A<�T�,�,`����MŢ��L�(K�	������%Q�����g�d�3o}��l���&V��T'�;^��'u�P"j�n9;p�9vw�s[ư�O�d����ħ{(��L����}s������e�@�yx>�[ק���V�]�ۗ�Q����N����%��e�eS��ϱ+�3*^dJ��*#��\8UO�GU��ښ^�oJ��M\^%�#�T�SV���TZ�>�te�'ր�u�7��tb+i�C���{�:!}z�P3�@) ���,���wU�^;|"��r��;9D���c�I&_F�ϭ2q��#���u8�Sx%��Uk͐߀�"0)�Q�����+����|���&>�x�gM����?�CG.����>�u�nІZ�A2ڊ�vu�V��a�U�9j��}엥���J.	�a�)��]I�B���s -����ks�S�Ql�><��ym>��!�x��
B3ߋ�R���(����~�	A90m*G��e*p`��WJ
��lnv}7���u]�:ؕw삩+Q��*@]~1�}�-w5ӹ��;��̪%�{��5����~u1����Yx�(E�۽f���!���K7����Q���Gc�? �"%���]��Ww|((Я�e�S�����.M��Fca������熹o@�f� `�q�e��Zj%-����i���� �C�W<�i MȎ�"o�?A�fʠ;�n��0{���o�W({�z���_�[�}e<x�]W��@���F��e��Y� z�2�'*��<O�-���G<HS|�˴������BJ���Q�|o*��t'k��Oc�miCI~L�J���Z/����TQu,3���i���r�D�"�A?j촚��D|g��H�gnᐊX}��jx��!d�(�zY@7b01*�Y�{Ǚ�T�X	U�_�̮<t!���2�en:j�y/��4�{�'�s�+��4�ӥ���Bu|ݷ/!\�!U���H���H�2ѥ$�
�a��Fp�2�F�q ���z_�uB./�P� ���x��7�TR�--���n�Q=s�F
�[ЃY��V���u"�!�ȅ!(���R��䦈��Q}�]�Iu�W� ����cM[wO�T�I7S�V)dP��7f�]Mx���F|�  ��	M�����JL�90哩K"(��g�ǽ��%������վ��k�R�c�A�\��O��fj���Z,���G���u�F2�XqX�Wh=��x��c1 �l��5@X�"U��K�g��̌I�b��VO@��B��t<Ԉ�dd��Z�,���E���)f���vڑ*�6���X� ���C�<��G��D4�HDf{�P�X"��\?ܒ��L~]_+ 9��B�]����s��Sv�'
�t��1��G��;"�'�$���+g2;3�y[?�R�Hf2����7a��?$���Y�.�&��ܫ�lq�(�P���.����@̇c9�0ZV���Y^�Pq��k�Fs��>�]��7�����H";�]MVI�;t�n�lN��Bl�Pݠ4t<.��Z4I��i���-bP�j6�
]I9�pVo��L�,ί��l3�'�ęw�+��Ec��I���oE�C)��̘{50p�3Aj��	�6i�8�S3����i[U �ދjNCKY�?s�,*�L'�|G�S(6��j�jW��xe����/s7?�&h>��$�� {Њ˘�n#�p�"c�ǅ�K����O�Q��)?c7V�&E����9��~��u���ּ�u���Ȉ#�� .��m�R�RfH�Q�ΔD�����rAR���8���4؜MI���g�3Z�	2�A����r�y�Ú���F�Ūㆳ\Z��[˿������k�(��@&/��N�|��L��<��P���Tx����V�[�E��&�C���b��1 2�W�w���f���9೥^Eʱ��jd8��d��C�R26��/4����#��L|��GJ��%=^��]��
���wt�f��bvs��9�����G]�C���`�i��A�p�B�m�Y���-��^s�D�*C�4��d�Cd�� �<�c�ЉKS����E�:�y�sm�Kuf���;2mN��%�ǘ�}o� -�q�!��g?3���?U7�_�=\�ߝ#ҍj�u�CS[��x����^S��.J	����׏�����ѕ�� �._��i�g[�a���AhX�f[4F����r��u���.��G�ְ��}8P����}#g�m�@%gq���}m�J�n�@�=�}i���gb��b�T�p�[;x�?S�&��e̎���<tl���a���
/I� gu�v�,Ż�����%��j���V6�ex�H�J�����s!	�J��g{��_�5#ku���<��!NU�f-�I�`|��j8�l�/�4_re�B΢��E.:�u(jȓ</6�
���؋u*e.U�נ�knG��8�ߏ ��(��Sx[""�6�s�P��w���ۧ�^UnKBT=����L��'��f5��Y�h�x�d��w��J�HöQv��'�l3cXHr/�G�E���-���I�T:Ρ]��DG|��ǀ�:-ږ�2^�5��X#�'��&jNB�S��H����WH�CS��ʟ{��������+b�;��)C���ԅ�I������bg�����,p�u���fi����)�{���e��`p�D+2�xB�>5�"�����S~�o:~��5�}"?��u��u�1�0�c��5��z��.ɋu�{���
���#p���`�D	�!_k���+,0�gf�ո�_���Ա�=��=B�?���B���X*���=��JW�ER�x]�!n]�!�����F�#&4��S,���x6�q���z���ΐ�Ǟ�u.P�7�`�A�W��S:p�1cF~7�h_�j�&�b��[� �PՓ��b�����i�eE��ļ
���7Ӻ�U���	Q׼�y���l`'�xB��)���ױ>��6B�<��;K#ۜ(M~,��p~�+�^o�]�ˌ��ut{Qw��J��-:��'����A�g����훃6�VZ2��焊��F�����!Ãc��K�	ueoz��ll�K����;��z�����n��}��Y�n=�JC��~M��S�$�?���]VR��6��l���H����Ь�G��y�ѓ�����8P�ڛb{���x��NTE�Lz�:r���461��R�H޿��^�b�r����W��y�F `LvǨ�B��Vh8Uw�O�W����8�񡸃�B��̿��%�殀�U�M�,�NS�1�!iD��aR�8�J��! �;�a�u�.]���(��4趁���I�`N;�{��0���?t}���������]��`ی*�4��6YT���4�q3�&��G�b����5��z"��C�]]eg�ߒ&�+�2�t�샚������t&����8n���a��#!����J�����&*�W�����"
�C��d?+5�-�Іw�N@R�ڢA�y�1ۍ�YǙO	�'T���9�]�A��B��>R�י�Sч����7ͣ�B�M9&��j<�,p�o`����b�4�����:�智ayl!|T�.�����h8qu��㝦۞i�[Uy��R�t�@�׀+3a��h0�9ֻfJO[�^}sʅ�E>�0I�x�~!@f���|l}�y1�Pݮ��"�^��p3E��%�?�h<�����c�d�'��5L�hT}����2��Z���qE8�n��X�jq"�t^eއk\ʇ{��\|�H#|��\})����'�^�D�6'S�ٳ�{Ϊ�[��m��mM�@(�S�R����[�����r��/��]ÕV�����ZQ�����j��T0$�@0�%:��zд&)���c���D�˦�����.K��rP�
�t
�����`Bʡ�Cʵ�Y�/M��B�h������v�@�'���1��opc5�C���ZK�K�7�q��4��1H>=q��N[�GXh�=bw��$��X\ڃ����,�F����h��پ�X�>5���ٺ�aۍΗ��:ӑ���AY����WM��-��ɅꝐOZ ��z��D#Rw4�gh��;(\������$6��p�'�d��(����j���q7�A�^�ǇA@����I�9A��$l���[�aºPy�/�������&�ד�V��˘�ڍo������O�>{����$�����nK����O�).H��Ű�˰v|+��?r.[C�/���vR:�H��ʭ���CW:j���~{Q'�|�Y~� ��憰���U��5C��e�g.�<�)yS����,o�D��( �H/WNY���E�CM�f��L�����,��i�5W'��d���`�O|=>��˼)�(i�8bKXUg'd�)a3��.?��Lj4e�s/�3���������%0"�e�ۼ�]�Y����%���j�S�4��_�ϰ�b/�)�2�Qc�m�ЇÊ�Ȕn�(���u&�*���2.�J���<f`P�?�� .P��tR���Dd��8S�#�J ×7�~�*�]�y�
i?�}�:]����)\���U�9&;�P�����)��v���_Z@H�G��4����
;����n���#�*�Ƕ:�Ӭ^�~��tRS�ZlO�cQ�|���X���H��n����Hh��d��5&
K-���!��1|"d>N��� +c؍�o~�I�#�2Xp��"!��.�}��nB��,�
m���k@TYo
\A5ʞ}���;bGI�xO*��׺���.�)���luM(b���܍��>�5��Bf�֭E�X�sT�x��E�W{�T`�Ț��-y�����d�N�ͤ-v6���Ë;w$\4xm�CX�g;���o81�N5H���j=�i�(���G��+r��B�.��:
lu��F�qJ>�2���.�>��@űdpKI=�A(�w\h�Ц������x�n2QV�����%I��e ry{� ��x�b�y��k�΋�ⶶr�t������CqP��G��F|6LVø�g�"�ˋ��?y�z��҇�Tآ�>��W:Zac������m��*�ױ�<��J��vT��R�y0�f��ߋ7+ګs������'�y�HS*�_i�N!@�Ҫ�m������;���8�r+e��^a���S��^5�F���g�g��.@��҃���9FX��FS3��-�7�<pv�`����<���I������B��+��7 `��2�[֫�=�DQ�|�y��%V�Wy�e3S�H���� וƗX-Lyx��4�/N͖��QV*sn�ER�١gTM5i�L��#*��⒴_�S�8��89- �kkK���w9�- �K{��2����6�@=Je��L���uj^�P
d�KZ5S�Bk��!�[�l�g�B�S���I��9Q����� ��b<��5�EwJ�k��MG�i[�i�B*�1 )���4J��\H����7V�ޓ9O�C�<��Grn`���u^���%��Ҷ\_�8�B<_L�]W��g�%���X�[` |����}g�w��R���_)<t�䊒���̤�bT�&��YQ��V��8��t5���28��ij������5��<��:��"b�6��c�����9���d������/2Y�&��\��ls�F/=������A�W����<�-�Q��;��E"�G�ۅ�@�4���ǜ��%2���{�5�Pnf�f����?G6��1�O��b3E��f�z�d�%V�P����mTn�PfbUE�B�XV`�͋Kr��S��7�E.L�@wF�7���HF٠�߼o-	@(�ܨ�ވ��o!�-�S��l��}�ڨ�i�AM����@7�s�"=�?*?2x�KM7��I�1t)��u�aZ�qt�	�u�L3S��qjͬG���EH\��jhi�8�s���

D�`��-z�e>h2�/���g%~\g�9��]
�=C�k5�I��K��_�#���EQ����&���%��U�%HU�k�B<.Y�ޛ:�-�Wb��n�	�©�R��{,�dp�ٗg�}(���A1�+8C(^�57o�J�5t�<,�S���S1�U��Pp�u����Ef����d���eϳ��%��|ǵ5�
7�쾖��錖�+ �o�cju2�(�62B»��]���֋�6��zP�� ��ށ|cü�R��{�������X�ڡu'^RE��m0��!/�Uc� Mo+/)3�m����`�R~
6��[ax��E���v|���<��.��C����D�ؔ�|�Ѭ�z��7�uD�=|tN_4�5�ٝ�5�K�%������J�y$�B�H�wʚ�8{���x�F�kA�l\��=kqH7ƪ�û��V8�%�*�׺'������r+|y���;�a���X�E��O��&f�@J�8g���U @���\�2�W�v���0R1�s.c��:�b�s�C���,ib~'�'Sh���8[�x
�E1�F������� ϱ5K��|�����f�k�o���>�[���8�7��[&�N<�x��ǫ7��a�w���O;����E��.�'��Tb�D;I�����q��U�_�����s���mGw�����Ha�STG��ƾ��������#��Y-�ϿV���fx�C�qW7F��M��ܢ8��������{�ؒJ���J	G�Ɏ��3K�7s\Uqn��N&��N���c9̗���_�����[o����#��ö����ư�QDP�?�������	9~F2�=��f �R>�YN�-��޳䫜f�TE]�tO̖��K1�{_"�(}��>�H�Z�����C�OAQ��[/0tV��dZ;gb���N��'4|�ΟM7��nYw�VK|Ep�n"x����
2�$��*�Ý�lt��/�1�����ר������������Ʉ���AX�ޤdoE��3���˔�.��ӭ�d���m��Kl��OOB�V����P��?����$��%�I�{}�Nc�jeD��j6���V4{�S�c	�F6��T���}Ri��7����_�>|�6��AU�@������f�n"��J7�g9@�)eb�n���݃��ε�P=W��"E�az���Rg!p/Ť'b�#q�q��1�+���b�-�.<5���;Q��װ��]��S~�r��4~Pp�b�ޘ'�7ya���|��Np0!�v\�'�<���Z���t�J�^�q�_��t�`]V5��ej�EA	��xWD-���E>��DaV|��:����;�ߚ[��P�l¥�ʾ��e�B`����\�՟W���R*R��	�Psh]�g���%��TǶ���O�?G��A_�^ՈV��<^��TaAq��� =�M�G�h�5�����ZQ��N�����}�B��[�%l�0��o�(Y�+��JL�
� U���
�guW�TI?e��/�FN3�gl�z���tb ������MiM���ۍ����qR�dgy�z���3�d!���2ʮ.@��[�k|ϼİ���g]!�~��bP�� �odOH�r����
�6��8�Ͷ��]��9� +ڪa�I�w��گ�Q�+��7u'���7�93�7�
w�1�jp?:�ճ�y�``���M�%�쿂vv�%��ZJ���^$Y'�7�T�ZkG��`�.��^��w]�R_�w��XcX��+@��L�_��PS�F������O��1SOؔ��k~��5ȇ��-�����#i�� ���i��@o_=%�0�``1iD>��t����'�CE�N��*/�(�y�����0*�N{��AY�&��Oi*�'Y7�!����M+<�&ݫ�Ұ6����ߓ&QN@"���U(.&u(����칧�q�ġ� 7�Y3 x�\&�񭋓�DQ-Ь��-L �)�I����OX�F�Fl1jh�w��(.u��%���.�Y��;s۸b�1�N�́�[:h���Ý4�z�cu߁��2�^Vsj6'S��"2
�rk�8w�[톗��4��.🌼j�'����o�d}MWe_I�6��gm�*zdJPq\��^�/���q¸<��
� G�n]Ǣ/'^���Tp��F�@�L7�k�3�I�3�w�DC���My`�_�G}�2�5)$_C�5�4���06�����-l֘ǌOk��x�6�A��|��Q8{K;�XO�!�Y�T:�.�ev��q��9�M��+խ	�:O��?��a��=�v�T®Jt�6Y�J�js[�,�<n��r�_���>�36-<�74T�D�=;b!D�*x�®����Ѝ�A؊M��մ@^0��#����|[i���;	��������5[�Gl`�����~g�U�*�ǖ�#Q�$*t�	r�&���8�>�$I�ڗ�^.V1�WB�w�`��������p��� f(��j�\���J��6~ N��^�~�#��A���m�
�Y�:6��]����DQ]H�ž��P�����*{P�~cB�"o���{�$�ń�lG�*��)"�!��- ��̸���)��
�`bw�?�|R�|s4���(��(���׹k����'.:0�1�v���g��&��S�yUe�s���}�>ehu�S��V^Z��x<x�1DG��}�&�j�|���bJC�O*���(���a� �����3�`�4����ҞOWϫ�±<��� pk([�&~W��֘m)���n�"t�3��Y���%ȱ*�?e���,c<�,b�I9��3Q��Q��1I�6=-��Ц��ߊ��upRz��9ùBs��*���&Z0�x��V�3.	%�"rs�r4P\�5B$A��&�@p���m������HeT��f7��C�Ͳ�_��b5<�N���39�&�0{�R$0s�Khw����s��T��F݄�	|���	s����i�;w�ɇ�R���,�����2���^/���Uю����$x<b�����^A�Ӟ??�*-ʋ���q�ff*��<�{��T���~���V�_�����k�1����X>�w0_��4φ{�
���N��8�'��5Z����PYƅ0V��n��T�<<_���On�W�2��n<�MK�.�� ����2�#�W?2Oh6]���;�D.�L�[��;�e��*�mCoٔ^g��	����a�>�e&ك��L��濯��0T���
��/���պ�-�$�9����OE1�w��mB����Jq���QÞb����a&��aB�^G���א����N�����%U�Ê��i°b�u���A!����9�5q��?Km���l��)��<陮U���ð�%�#@��I��R�ܼ���L�V����{jeV�O��i:�*E2��+�o�>�c�������P�Φ}��q5��d;���caSD�P�+�N� Gb�4K0\9�O3����2�wd�I���3N6�-*o�*s�Ӝ<�=�)���	`�L\�9�QC��, �1��Ծ�Z .���t�c�a-|Kau�2��n8[��6�X3�}v����E���V�]�Ӂ�ڐ�fQg��%�"Z.���q��ڭ5��[��uo%��3:z������p�T�z�1�0{�Iv�,��L�m��x�$^��T�u�̜�c����I�_8灂�-��]�����>nƷ�$A��h�w-��r��z[�a�=��w��"�)���GT��r��N {��ۋW����d�-ѯ�޾�f�.<�>[s��I��a��v{E89�� 0B�[��s�z�K�k%��pSS��n�,�u^TP5����H������h��4��3��6�l�*Vc�}�B�S�4�/����6Y�`�Ұ���R7�O�u�F;7}hC���ڍ{YU��XX�����0{[QSa?�mnѳ�Q%F�?�u��\�U��_�ȾiO���F��6�_DpI��������R̦�L���l��j#�A��C��6�_6k�s��=bR��y���eW}�����.J3���׭y����OQ��VW�5H��D<��^�<
����*+O��P���?I��)�丬XEh�)LBG�>hr{&w᠜�1�)��e\�ʤ$�_�ㅀ���L&׼!�;����W�
QU52�A ���N֬I,�%Z��1��y����p����C�3�z���NR��g�תtG�� �:�J%t$�n������ĂW�Q��(��GUv�DVվE�ՈR�ώ)F�f.Tv|ܵb�L���´�$��Q��_��N��9�Pb�@3_��W�@��g��� ���~=K��J��'t�ِ���{+����x�A�D���2Q�-�;Y��۬�Q�g���ǦQl�MT�!j���| �R3<{�m��h��6��Q��A��=�dTbp�uz�q03j{S��!W����U�J�B��u���|jQ�Z,����� �q���r\Zd�T\^ss���p7F�K�?"#!+�
j4˪�H"B�~�'J����N�b$C�
?~��4r�������[�)L���ķ�h�Bĺh^���s�-�����\b�]A�����y�Lɫ�K@`�G����Q!v�G�*�"��ەp5�`'B��@�jgau�������uRD�K��?�!��v�U�p�QD�<g�f��c1C"*��C\�[v�?,����Уמ�|�fKG9d?��y�ި���X�r�)S$/��!��E��D�'m�Oyw��M��@��4~�vq-\^=o��D�J��ۛ1�"y_��Q)ي��.�tǵR�FL�pk����>���JD�BW�O�^�ֺ4mR7�	#���C9�t?5����`gF��a0�	֮~�Pri˫lA�s�G�[G�R:8N����W��%���)�A����"Ahs1護�r���Q�:tM�/����R��N��� K�������aɂ�Q�M�T�=���� I�`h<櫉7�b�Dp�B� ,�*yG�j���;/GE�~t�[0��PJ	��j
9_߾F�9�|��g�F?�>��ٗ��c�W�ntS�qx9%���j!
}_�z �8�Q`�yL���hy������Q*���X�R�wx�߁��i��d׿�Z�+OX ̀��~��
�i�m���9�a���̇c�����V|/�c��H~/�������[ ��xub�-�L�]P5@�4�Y 	@�D�3����A���2+�d3����Ge��`c������ŬE,uLӻ�^=_Ξ��椩 ���Q������%hj]�3���K}E�W⍽ͧ�	o-�8�B"e�)�|��^����ڑ@�!ۅ��W��o�`�	�<n]�>#/��n�pc�և ���A$���>��d|
?�j����f���v�IB�1̘)���}��ɰ�[p�iC���nQQ�Ք��>=k=A�,�W�⧇��Q�sIvZd�ڷ�m����M��Ӫ3\�ڇ]�L&H����=��`��	�S���1�i[�RO�����YE�\hL��$?�$#��S�G:4K����G�v�O�E�1:*���x�.FZ��l�0��N$�����H�'��'?��*.�	�`���D�\<�w!��0�)��F[�Vi�(H�>kmDǏ8M�U�-���7��qfj�O��*u�/�n
D��SSˊ����X��}&�Z��]�+��f��=[�	�ךw�49���>a\OD� �V�<q��hdD"o�P*@��P�}' �}-������+���a���#?c���,��1Z��b(�������5����>��J�*s��g^NB�c,��.���X��{	Ȕ�[}d��D�5�����`�������7G[6�}o.�Q�H���x}���I>�s�7�؋t����xP������X.����;��E�/��������qUi6��jMr�h`\,�m�ޖd�kG�b�wc��T��̝��O��27aE��׶���m�!֍ұ���q2ӻ�~�ù!Ƕ)z	�ͺ?�Wޏj��e�_g���Y�!o%�d��SAr���<y��
U��5E�`]{i�q�]Ux�	�'�ѣ�4�ݗ� �D�+�¤��%�@�"�f#qZ�51��7�P�`�_�T�KI�/͝t^/=��<.�xNN�<��]|�2N��ȡ>��]�01�j��f�RZ+�2�7�J6(����ҥ��}R/)�E��E�r���gǾ��h�t����&����o˟w��v*�x��;p��}p�46(ZQ���7���H�BgK�r0TX�+3��?��V�?g��c@�%���'+�u%_;�u����K��Q(X�H���Sgi�}ib��@��C{���şC3�pr�So�Ӓ��!�7�I��%��J'���u��������;�+�v���{2Ux��+�!	��B�N'�ط��*��:BY�:�S�NU2��5��:�J#�l#�B,o�����⃚H>o.��W!������'����:�Z�>��ׅ&p��Ov�ħC����q��Ч�)��nf�Y�6��At	h=i�b��NɕW�5����d��E��	��I�F`�����4z�u��j]s��M�o���lL����.�x'Z�Ux7��������l��|�C�|���o.?�z�����b�.X��ٓq\A�Ƥ�+M#S�O��5)ӈa�e�xAhT.K��	a~����ap"�}�1aP�$��۫Z��2�,����2�F��,I\n
�5=1e��w����Q�U,Q��#�5��B^<��V��?�0��	�\r4r���^�D��=h>�[����b'���/�)2IT�P�%!�,���o�xuMy�"�����z���x"Iѡ--�k�	3��
�]<>b��9K3YnO_��wі�>����5���Ha�{�k���o�3RH�pe��U�&9�R!7����<^�[���sέ\�&�	��6����|�`�s���Jf`�0`n�&���/y�.��[�_莜O�R�l��_e�@�����>�}�J+�i�������.N��*��Y�_k�E�Ɍ�k�D@�{ⴁ�m���~�}�*�&h��2��[0&�4!]��=7��4u��l�&V�+ӕ9%��P��|e��Z�|+Y ��D'�P��Sx�e!����ʗ��H�0�K����q�#zA��W�����W�RG�:4��m�]���EvU2&Ԃ?�<Ď%�%��8�N8�;�@�,-3-����|qc�B*���ů�J�*���["=\�óWd�yyV�:M\Y�b���hӏ]��>����԰�2�ak����{����:p�PJ��6�%�H��M
C��͢���ŝ���y��BUE�����2X
����D��ͯ$�'������]��2���z-8W�܎Eϔ����;����s�l�PG��D�ь�O���9<�M�^�Q�\����v�S��&�I�u�LA�0�� kէB�;Hv����9��9�hi�Le�����'b2g�R/8��\�q���)��ם�Fu���ݩ,��J�3�htN(��5�o7*��Y?�q� ��ǹc�w!r�2���}����b��L4w���2�0�y���e4S��HڿÈŚ���S�m&	�\u��xJ�5e�Li�����A�ĝ@�@�b�H��9?h�nh�T�&�t��	?$�ů�h
r�c�Jkf8��_���7��y��i����!�2t-#�׭��hG6��@��JI�����D��o���	,C��-?�M�ըN��3�n'�؊��V=g�N܂c�۠۷��B1ѝ ���X����چ��
�Q�P�{