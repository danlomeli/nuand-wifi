��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� rā�SZ )����C.��&0C]�-��[�3�-���+��պݣ�k�J�vo`�A�����f����u�X���v�=�а���]Q�Wۿ�߸�=_Q�X����j>��Zw�K��SvX��ƥ.���#�����Z�0���#7{��\S$��@1I�QX~TQ�E��db����۰� ���>0�%�9�j汈��}��1� ��2���h�G��SeY�a���	'<x�p��k�H`�H�j^y�0�s�78+���ֳ�`�R3dW��_��{p[�?$�s0��#�zS�_��bH
�c�p�IL7]� |����Q�� ��Rr���=��E즕2%�����`�^��l�q-�]�p��jf��Ӽ-f%H���ȳ�>��+���M�71��4_�) 3�46h�rb�J�W� k�h~K0�>P$�_n)���5�r�j��W�J&޴o��$>��6��ŀ�;A~<6P��K�~��f��*I
�Z��}`q���ApC��n���g���3��-�іrO�mF���,�$��@�BI�q�}��Ȥ֐����î�䂧��@������U���vU������ �T#K@f�㯁����|95<@���+�-�)�����K���FI�k���*@�m&���
���ma1[�2�u�I�\�U�yu���o�|��2����;�W�W�}P�K>%5�'�8���׫=����k��,�t�M�0�8]q3���N���GvZ�i�+ C�e
��Ќ�S�v<%���q��e_��
�k�夞��>ZO7E~��5k�TW Aod��eE���G���ɑ-'���?�G$����ќ����8ɸ+ 5ʗ���l�d��,�J�
�^�3b,�����J����#n�zK����z�&��;|�\�^���'e�W�����">�w*	FO�Δ��v���I�h�*�hF�������	���B7��c�ppĽ^� �W��#�2��t#��w�ET�g$zM�%��T������( ����zwӶ�f)�Ր�-�;T�d-LY���`��B5_��%����<V�{Q��y����������0>"m�B�f�2�"�8���Ռ�2��m � D��v�@o��EE�>L<t^��!~g]D��b#�0�GxvoH�SuJ�V*��8{���K2�W�i�9s��="��o�:S�u�HN^�4v�΃������4���3���x"�����l�4�QqUqؙx��F�C:.I�	�jXX���������E��2�L�s�%߇���"�LO��l�}4�d�ڨ_�����q����6���B{ ��4�%<�S�h�����Q��������T��RLJl{�đ�+���!%��Q�~lM���4�����@a���j}g䉅�A]R�X4ɐE����[R�~�Y��N�����<���o�6S����$���ζL}�ɛ��#�u�1*&���I�"1����)����Иβ��Q�����j�&�_U�����}�-��#U�b�׫�7��>����P��G�y����*-z��h�d��'˱�K1{I�%�a�ѥ�=+l���v{
��!��t$X �v��I�����)kV��;�={�;<A�q��	C�\|�w���ݬ�_��?'�4�]Wr_��+���CZ�$�)���|�#�+���fk����[۔�[#���7��<�,3�Fb��&�w�����ݵ�G�͏ILP��:B�r�#N?8�$���KPv��⺐kQ���"�qU�IK���>��!>	()�v��O�61M@)�j�ua��`�4h&*�ǂ��|Ymό-t�?m��	5�#DAk g|�SgT���͐���*��G4j� ���M�����+:�VN��ԆL�?��c*5�S;��,�o�u��S{��ޗ!8����&F� ��U��.�'+l��!g!��v>>n8� �����.p�O�'��}�� w��;N��?��h�;��4�J>��b��_]�q�����E�ǔS0ڒ�Q0���� q�e��q�l�6}�8}��z�����Ԅ�Z3[�~����0Rn�oL�}C?Ob�����S~�&8c%&+�[D0Z�Q���7>����I�YFj��!r���m�[P$]�(5��ޔx�~��n��풼]z4M�2��W\e�)#<n��M���j�Γ&,���M�����I��ņ{����\�㓺�	�t�a~֚��<�E)5�GJ�+�pn �R�����L��E��P��ۻ����.s+���S)�U��z]��-�w�M���M[��0��iE�<�LC5�0"ڟX!�ԩ킵U 2d�V%��dJ�G���GF���2u �/6S�1�J�.p�h�Is�~�b����R�V�̧U�Ŗ��}����Z'ܫ�����C���C�G�8�ѥ�*�t%V����I��˱c3D�����M��r5�*G�A� ~l6r�o��i�`�pl�t�tj�""�g�A�+\4.�h-���Ek�L�}񾀸i�T4��E�a\`َ,걂�,����R��&����f(u��p��`�(c$z�nk	x��Ø1/|�d�e� ���)���y��L��R�1����{��I�rD���o@�# Nxf�a��]v�
%6�ț3�ܕ��#_���N�4��W��9D�Ymk��Y;g=S�X��C��L�ޭOGUW7�6_����d�=hf�o�f\��D���b�E�iR�a糚<#<�mh��U�Q�O�O��w�s.���4_��X�e~ؐ1�b>����wl���S}Q�3;�:J�gGӧ���� �/�ÍՔ��Lr܋�{�M� aF��mG��U��1�W��R�3�~���ߧeQ��h/�Ѥ^�y�:XL�S��uȑ�)_Y��leP� 0��MF�(vΒ9p��9��O�R�E�z�oj�%��\W*�B\���&����ַl>~�EI��s�3WxU�=!��&#�f�8�P㠸�+����c%�sEk�1J����k�ck��3�b���v���x��>��u��}����/Yg���H��چ+��;=�l0���8��3-N1r�s�z��?�[�U­m׿[�eT�%f�Y�X.QVM7����]]����z�޷����K@����9!<r���"j������'��A�=W��p��tg:U抷dX��!t��s�`�Ooww ID	:���;�hlE�o�1�o�l��Ę���A�$�d��|G�T�` ����ql��'��Ɩm�1BǊ����.{�mR
Dv��yDp�9lL{JT�<u�F���xiJK)y?XDQ�)MT$'�TJ�t��f �]g�h@o������zU��;���&��a0�?I���?!>��?V���}�GTє���^���{/7��A��ɔ"�r�1�&�:c�+��;Y��%���?�Vh�0M�֭�vu��pe�:�&���b�:V��0��v\�g��!�+c~����oVҢd��U�h�BDP�k�)�s��(l.(��6�Q ��$W��-�d��yO �3)%Q�L�	[�/�l/=��q�����2#�g��Ĭ>Hˡa�u�k+�o�Ͱ�?N6�	*b�f�k��#��ƣ�F��x^�2B��^�L�kn��sD%vB��4�Y�`��D��`�BT�;����l��Xț�T��]��C�����U
��(�S��âf[�(Ӳ��|͡9Q���,�i���k%��ֻ�G�H�$��ٻ[���pq!?O�(o����]���l��m�r>f/��u�\�&S�����2�����-��$�d �]��ĚY�J�Bu艠�Ώ�q��4$ ���bG�T��}����o�uv��<����V��A����v��P���4�l�c{��aD
['����Z��'w���՟����*s�ji�Q>�i���mbF�3%�������d�$Ϡ�����
Z�����x�w���eH�<��#[��N#uyr6��`[r���������-!���x&�k�-e�ᙼsh�.3�):��׈3e.3��m�m�UWLۖx w����o18�)��F����X�mO�1�}�/�v�X�(Ώ������T[ �S�w�6��S�Ul�yq ��Pq%�szD��t����٠.*%���|��q�7���⿭Z��0<�x	wy.Ξ��X��GEu�E����0BG������(k�Ҁ���x׾�E�Q������S!���2;aݜ[�����s���D��<,�aj7��]E3���4Wa�Υ��8�l����=7��^�%	9+{�T���n"������3���Ⱥ�������Fg��'m��i�v�Q��������+��]hTk�J����AZ��2E�Ng��$3%u���Lsh��@����0pg��^��P�x�6���1���l�bl#��5��შ#c�� �6^���$�-��#��vy�Ċ�(I���xNL9��o`al�~����X!꺳�������	��7+��-�>J܍�Ў���/�ye���4��CH�=����%����N~8�)��B	�=;��SU-V�׵�b� ��9 D�O4�7�o��3��_���I��I;�����$LF��\����l<x"dO�MG	m&ͧjN`=8P������	ex���X������{H�q�ՙ�n5���xL��~��H�"7��YOve?%r-��j	h�Q`��XR3�_��s�v���ʼh��2۷�DHW��	�u*ͻ�L���[o��իX�D��,8d{ ���<V(v�e�D����v�S�	�j:��xAx���#�\T�(V�lY:/�|�ۥR��Z)u}_�g�8i�b^u5�u�~�Kc<��:�
�au��!���x]J��s���K	dQ�x�wH�%��o���A�7%Ư�~[���Y�x"���QxFʐ�48��#BR��j�V�Q�3螋�c��(֣�7�.�2B�(�3�[b��e�*����
c֖|c��G|��L Ow|3�����X<Y�ż I+�\������'<s@q�Aƈ�N�+���d�"e�XrFY�W�FӜ8B�2:��ʈ��HT�
$���=��lN����տ���y� ����2��:�n�{4�ѵ]�A� ao�K�\�"�� �h�Va��?���в$9��/p�	�υ$�����K�7�`pU�]���jqz]������T��B��-�����X�+����t����f���3}_{M#@6�����p?�X�2��j;��ɛ�2V��5�Ҟ7�a�KQj��Ȉ��Ӵ_\C5�O�G�J�eP��M:+j���k�,��g��Q~�,�D���T�� Ùu�D����ZiPBLR �]Cm'�=r�V^���E�i��1�R���K�g`/��e��w��A��^<'z�5%�p�����Ȼ�f�"�U�<�;�/�7�<�r�(_U�l�l�7j���0��a�OQ�,q�~S���6��kYK.�c/Jg�hNE~����� �L�I8���eЬ�˒�}d��oL��{�� wg{9>� �#iN�&pQ��x��;��Vy/�`/�wo��9��c���Ʌ	�sa�i���b�Qoh��ϑ�U���qю5m���k�z}Im���E9�^q��=�Y�Kۇ,��i��5�cy@Ί>�:1�_b_і���k����v�!���[o��zĦ?�Q%>�y,V�MsG�*:H�#	���W*�c�m�
�K�b��Y��YG!���mY$����!0�?`,�����\�8�F�֧x :��)�րy���7U$Spt7�8�Y�Y1�9���J��M�˾+�
k�����ޝ����2.�_�����pWQ��T*��<�Xl��A�P}�#צ꡿�@�P��g*?���j4Mpw7����� ��G�&Oa� XW#��u���#4���|�؈�/�筳��t���6�-](v|�Y�8_��7<R�3�Q��i�f���bl7u'�����<uX�%�CFZ �Ofkw���H�J��j�:�=��P�����v�;��a#g���ҹ��x��i���-�{V+���c�(P��c62j�߲P�d��Q8�\)ox$��~P��
t��Fl:�J��$?�U?���>��ۗ�eaR`�HXS�K��vWE�q߅:�#$V�f0�0����#�	\�BH'`^�.C�x�{�;�����C&��̋�zC���659��1�G��c�π_о��~]iw�����/�W�R��<up��"Qg_��	�����x&�E��>'�<�m}�A��{V���}�ʥ:,`F�O��nA�4��=a��2�E�1�(r���-��S�s�y~����E���g�F�&H�#��	��z}S�̒���� �+���芊䛭���{�Yf3�Q�R(��9pP�~$`�P@ݵ�}�b��|�	�����ب�ą"��q8��i<���8����|"˃�$�V�ԭ�|��A�}�d:0��t�?��>��3u�O�9�dg��N��;���4�C����[���x�d��m�hN��Y�����C)�٦4��02�:9�T�/��)�.��)�"�Ip����t�?!����(�=�k����~wT�g�������"�Tt����`��J�+/]:�jz�IOJh�:�9�?n���Y ��`�g}�����B.��9���s�$G�4HjI��c�E#��|ߊA�(�6�⦖1�Lܒg�V�޽����2� JI��$��ڞ�~�p���c��������^/��j��Rʑ�G/��H8�S'Lr��1=���-�C�Q��A'����_���#��sEϗc�*KP���?!�?��{-$j�H`�_qͶn"-V�!�>/���o�&����?���SG�Or���|c���X����,�U�<(=�~s��n���}r~�G�"\7{A���Lb�#�3�`љ1���@?���[c��{��ڣ�;��'�9'�}[��ؐ�g��_��۪6e,l���Nlo�\K ��Ua�Hd��rh���@������u��B����Qw4?WPQ1�!�m��;Ne�/�-7�Nu��vUe���9xj/�Wj� ��>�`���f^
��.��Z�L��!�EK�R�x�����k�_bT�_�, �ɂ�Zپ�L�}�&pK��*���� g532ܵڵ�4B��+�vQ���vw��T	�yYXx�+��;L�������a�A������/��z��[�-�t��s��?���ذ��9˸��|��a��µ��Ep�NK^�g��`5����{�Nͤf+ʒ�V�ߚ�y����4���]���RZ8�\O96:�#j�����n�2w�xm��$��g0���m���<3�.p�~ym~� ��6L3B}��Q��p��E��^�C���iS'Y^�P�r�?G��]�Z<�Ǆ.ƌ�g��nɧ����U�{�s�r�O6���N��;x��(�C�Vc�VC���8��ԧo�M��_JbN ���]ġ"7���yT B��#��K5zf�����I8p)�W�3�d%�N��q��=aM �Sf��m/�C ���D,w.l���H9[Ҩ�Q�+�`#�x<@/�oL�A�vC��s�V��l`N�뷞{�� ��^ܩ}H�aD����BT1,]M	q�m]��c���DO����E�*g�ϧ��a7#���x����	�T�^��8��0��2	����b��-�&��	�/���7����\t�w��+�f��}P{mW��'ꥶ�يM,�@��9}K�]1����$����Q5R�&�_'4��|g#f�~�nc��� �R�\v9/�2VeFe/�:U�;JCv.<x�^8Z�:2�"����>>�AVa-�9n�a{���$�s�Y
�0��y7f����ɤ�fێDɱ�b/ܭ�I+�q؄�K��:�}� �g;F��7��h�����&�4ߙ`�ص�V��w.���Q��1E�z��ن��Ձ��O�R˶&.S���5ۖ���G�;q|+�(�@i�y�u��>I��Ō�|��ј��Zy����Ȧ*/B�v��\Y�Dv��J�C��Q�G�8B���@!l����f8b�)+�DSp� ٜAyM��3����n��˹�N%��a�I=��hw�S�s����o}�󆢓���k&a܌=���`�#������W��������ġ��a�(��c�o��`�8�}8�~R��>��/q);��Wp�0��f�H�`v�j�5>�S�so����w��S�9F�ƍ*�Հ
���w%M[�^֚�E2~-�w@�r^.�6�E�+�n������e��1��\���#mI�i����U���3����
#�I0��	��u*(��m�:+�`�ŸC��Ho�ע�C��aTK2������ºC�>[[YH�e���$�d��K|G�&Ȓ.a�������.EU֓�/��w�S���Z�ѯ����C1%�'��N�ĕ�91Yå����i�JI�$�3�dk�wuփ^�n�δ��¡�|��P��1��E���E,�A��Pm47= d���qsA�n����W�-=f��4�>�o�=���i�&��̃*e�"LT!�7+���a�Q�ȼЫ�q��n�R�<�i�_,f�N�I1��s]�{j�C��A��0|L*5���g���DxwG~G�:'�D�c��7��O����idNy7���.�;�=��#k�K�QZ�ˎg�l��w��Y����۸[!c�4`�������T�E�X#�@7��-RT�>�ȅ�`�S�6�"��;$�*�=+ZV���Iθɞ4�dF�"�C�bGTL�^yjT���p�@u:����-��������|�r0K�� IA�r��l])���|�;���$�G�Zz�]�;U:�`\�[m�����\��}�����#vHQ2T������M�A�M����r�]i�%�0KJ�kZ�ŵg Jzò������]�+����]FK���XflClEJ�y���y� xR��������b�&1&����[��1B�ߛ��	h�Y�������,�}�<���9�W-���>栬����E�oZ�3�@�v���{j�{=U1�sG��0+4��g��l�����du�3C�B�{���xFY���"IlT���M|Q���t!�T#�ݨMK�