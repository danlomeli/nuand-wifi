��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� rā�SZ )����C.��&0C]�-��[�3�-���+��պݣ�k�J�vo`�A�����f����u�X���v�=�а���]Q�Wۿ�߸�=_Q�X����j>��Zw�K��SvX��ƥ.���#�����Z�0���#7{��\S$��@1I�QX~TQ�E��db����۰� ���>0�%�9�j汈��}��1� ��2���h�G��SeY�a���	'<x�p��k�H`�H�j^y�0�s�78+���ֳ�`�R3dW��_��{p[�?$�s0��#�zS�_��bH
�c�p�IL7]� |����Q�� ��Rr���=��E즕2%�����`�^��l�q-�]�p��jf��Ӽ-f%H���ȳ�>��+���M�71��4_�) 3�46h�rb�J�W� k�h~K0�>P$�_n)���5�r�j��W�J&޴o��$>��6��ŀ�;A~<6P��K�~��f��*I
�Z��}`q���ApC��n���g���3��-�іrO�mF���,�$��@�BI�q�}��Ȥ֐����î�䂧��@������U���vU������ �T#K@f�㯁����|95<@���+�-�)�����K���FI�k���*@�m&���
���ma1[�2�u�I�\�U�yu���o�|��2����;�W�W�}P�K>%5�'�8���׫=����k��,�t�M�0�8]q3���N���GvZ�i�+ C�e
��Ќ�S�v<%���q��e_��
�k�夞��>ZO7E~��5k�TW Aod��eE�z��ߎ"c��vX..�wy4��VT;/�XN�p!.��e#\�����[Gi������dW�nT�!���O��I����ߠ_jvni`��t�L1�)�=��q~�[aDG�d�1�x�mPa��jG���O��x��ZL�M��٢��5�=����-'$��S�j<H	��Y�8A+o�]e[��3p�a9O8ޝkm�Fdl�|�r���c�@�ӎ9���{w�5����S����6���oB�`Z�e)o7��UN�ǫi1�"��ӕ�aO#�h=b���D�wO��*ש�Vƽ�g����h:����w��[� CV�����!r�Q��C~�=�^���`��3\-��ؑ�HG��y���
C���Y=Y;X-^e�*1�}:̘jBP}��ի�A�ؕ܏v���X��`[�9b+��p����r�u��ngz���uk�'�*�)�?�.~J�\f�����|�!u5t'��u<w����#VYqxB=9m�FJ���Im�qA��1��CmW�W�w:C-��ma��\��@xs4���GR� C�n�Q�����y�b���D�8��cD�m��*�?k�q;D�yC ?�6+�Sq��5���\���oaĕg�z���r=���D�Z NmSϽ��/E��ԏO�V�uY����y\�����M�^[�b�4Ʌ�M����\dd\�9��?�I��/X��ɬ��+>|��`*���$��{���9�:p��8nz2������rB�)M�\�S�t��`��R�}X���|>��t�T��U�	�O>�p��I_YT`H��9�y�V�:�R�����]Jȧ�m�YUg�=�٪K��Sh�!�ߨ�R��$ck��]>� 1�F�����HQ�ξ4�)>�Q��f�����L���dOϳ���r��R��D��%m����0�+$Xo@q~���"���/�K�����/�5wK�p��(����ş)����Akl�.[>�	��[`P�m��(o5��K��f�3V=8l���D�1}	M�W��
�M���,��(첝;��ҹ�K�-�0mo���tr��x����౎ɜH�J���W�l�c��Tx�c�"�Mu��ހ�[J0=~���5=h�f�7+�K�dH��N���y/����	1`��:lS>|��R:����m���g���AP��&�ox�1`�rSRv��**ѭ�F}���{�)2�ھ#2Va���[c�>
���+�PyrU=ׯ���y !s�{��T{�-��"���Y�ߒ+���k�<��M��He��l��˩����<�������_'w�7�*x�����n9�7.�}���Ȼx�=eZ��'��I�u�o��`$���f`����_�dk�d�'D��ɜ0���'�A��S-A*E^�k�7��3=6�_��S��:���≚S��S�1���M*���uy�=�Eew�kI�����5`��~���n���"��ݼ��u��$�����s�AO��ekO�
U��F�}@�￯̀��J��ޛ�2<�����y��q�ۅ���A#�1��ӱYN�n��ԉĢ��F�6��w�N^?��u4��m��}�J;�>�I@����&0LH#j{�"�)�%���Y��$��V.��FKM�;v`S�g�~���;�5�Px 	K�H��|��B�^�=����]���>#�Rp�WO�<W��V�md"0�9/�|ם3�;l��$�����׀��\X��=�b� �t�����o^�3y}�lkJC����q<��� �+�Y�5�a��k&�n�z�j}|ߤ�T���a}�������:�:k�GOB�}���7O7gA���az��u6��F5���c|�4�{:�ְ𣡓$�:^.bdǣ���1)�d�W�-��|��4=	̶�7Ud��� 9F�"��4'�ؖ?�v&`����������/��t�囃��fr,Tmt����r�y�ԉO�3MiO������H�y�O�n��{���E��L(��ڂ���4�j¦���T���M�ɩ?��1����m#.F(G׋jn�q���?���Z��v�-�wt��5����݉�?S�yC>��爜m�׽s��&�N�B�@N����!��<�K�:�?�I�5=�\���H?H?�p��b�'�G�f�����܏�.�<o�_o��ߛ?&�
ԩ�\�a�O	�ܛq���ȧM:�).<@�`��W�>�?;A���@��v9�M!�4������[,z|l;�dԌ�z���{^�"���ܟ���%�{uR��� �G��t�	��ڑ�U�h1 �&��Xw��a��K�0M����}܅�.WO�XG>�Iґi�<�P�:l}@���)�H]U�9�
��#(|u��s��x�1�.��L�bm؝�{M��)�>r�m��a�����Ce�X��S��$u|5E�-�s��iPV�F�^��_�auv�����L��+}m¡DQ�0ō�q���0�s�ZD�����I��b�Юj���9�	��wgMR�Ԫ�����A�K��F���9��j��f�C$`Fp1=`�
�i�δ�=��A�S4�f�$x��T8��<����V}���j����]�d���	�ވIь���[q���4���U`��!a���q����+��NpC��(���."��$���Bٕ5��C��sל4L��!�ؖ�3]�r�������0
1:����$˝����a�BH�O�c*�JPe�L��fw�/��b7�	�D��Pc(Ġ�DI��P@�ء�#]����H�w?{�tE�T]3�ׅ���J��y^7;�-�6�b�z�B��i��z����F�|�:�ft|лb�R	Z�?��D���z�"�h�f隁֡�'��7�Yd!I3C�~��/�(�NWLY?3 �&��yP�����8��U�V3O~ŝ+s�k�z�0D�c��z�l$��!c*���̫瞾NxpN�7�^-�ntaք+O�A�C�u=�(�	����7/^]����I��ր_C�kîtjd� �5��yij���N�5�,�Z��arfh%��!�8|R��y�`ʲm+�����L4���{��ܰ�����0O���G4�`�~g(-9��;H�,�(	<y�O����j��F�������`����壳�d;��я
�n����&H�˭���vʦL^J�!�6��1�/W�u�H����]����J�$*��c�鸦������` ���3��-o�1��b���>/V���(&L���|���E{��IZ�d���;����S1��y:�wv��>#9���:�;tm�}	���4Jwt��^��?�Ǧ�u���TL��n�W�!���>u��UbDg��hag���SK�h���o\#�ì����v�+���Ֆ�f!�aN~�2o�����@�(9K4�>{V��2a.n��*C|���ݹͬ���1Z�U�)~+�8
��뽤�%��!]�A�Hd�=�A������`�:��(�S���#?�iJ�?�N�8��	���5�k��Ј2̒�)�l\\�2�~F�F���_��|��D�q��7����)$�gݺ�z��\s1K�=*�"�){�\���A��� �Ϡwi@�c=P}�6��(�a�
��EA�_�H^1�)��Z�ᒶf^h�N���j����)ԨV��ӑQ�d�.��x�(�$�t��L)�	�E��B��,�ے��f���=ؓ}v+Ʉt7�"������2�q_��xKP��/-:��,�4���3�bb����B�#���Æ��&�B�N�̃�t�@x*զp�0��H���.%��#>�.. ����R�Խ�q]�%p.��hQ��!2SԲ�L���nm\K���MJ���{�N��08X�
�H�#����a�V��C��8sMő�őJ3�o
 ��������̣[p�g�:BĶwA}C��iu��y�t��P�ΟSf�f��}�)�E��/}A���?���vao��[t�]�[\��+��[M��2V��Ij�ؽo�Ȗiq��7mf����X��G��S�c�,Te�-ْ	x�%؆�?��b*E��33�/i%�mB�Q{�W܈E�׭�����P$�g���`���U�4�ȗn�v�Z�?Z��n�W}��� �r�� ֓���y'�B�Jv�03�ȹ��&6��h�0^_��4�Wc�L~�*.���:����%�	��QL�U�7E�L68���?2�/ǽ|s/.�CLi�������%��g������� )�?��_%#�F��n�Q��9��iTdYg��G3A7�X��)�����v�t:hh�*w3�{C��R�yP�	Lٴl	�1ڳq*��uJ��ˏ�(5�c��9��]]y�d�����&���i��Mg�~����6-��d�x�Z�vhjVP9�L�t/����J?�:|
hE�Lj~�q�B���g���M���Y�ּ�߃m}�Okd�˒���;�C�:���u4a������Ŵ�I� �%<�=�X���$ lWDMV�_�����c�^�.Q	�*��
]�G蜋�����"�iԨ�Ҟ�n�/#��z�y<h�F�G��aAb�����^3��U˲$����i6?��)�.kLOۋ�v��?��I�?�����z[�ҏ>5&�O�I�V�o_c��|R���I���T�d�Eͽʇ���f�*q�Lw�j�e*ZП�a��~`�?���ؐ�~��K|/��4�x�Bb��A�A���ӎV7z�ޑ�2#GtP.o2��OTd�V��$y�{گm;/b%<��Sc#CDL%���4u'<�p>����H��*>�09��:"�?{�׿�|��f��Nb�%yym��%f��U��
�,5�b��x�%2�O̼/2IBX�g�3�y�8y;��=E�g��v��bi�1~�	��n��ŐAd���
=9�/`Ď�?�ٰĽQee�X�i%�|�����rO<'�'β�5�6�~;(<~���e|Z����K��n���+��.j.b��M�,���u N�l����o�,��<#/J��A����DU���Y~e��iG���;k4�-#mf���G�Cm��G�/�D��4u	��=�EΖI�zՆ����^wt$bL�e��0C�T��vh���N��B`hڬ} ��n�>�̸(�87�^��g)���S��
g(�o��X�Rӛuҡ�6@��w�n �Q���I:`�F�/&at��Two�(�2V<�'�	�b���0���ɛ
�rϊ+0]��p��p.���;�յ���3{O���*�aY�FO��r�� 5�;˙7$�vy�3��k2@��ha_}��Y��p���$���+���~;ğ�(�+n�aͧ<�+4�pc����z�R�d^%�y��k��� K�ϭzZaeI�X7�sņ\2ˎ�m� �b��wwiFē�%��g�¦f�[��Z��5a���`���ew�^1��?9�0��=��� $�"�c|�S4�I�4%��?o�k�z�J#���ü����<$h=s�I��l�1	�V�΍�T�N2�a�����t�u� y�%��I����t��Y(�X�k��~��]҄p���4+�5w\��E��+X�
ϸ�,c�\���h����@+�ݬ�����Z�T3�-o��
���Q����t��<������M�[Kn ��4rV�1#���;��5�����D�X�ޖ,ux]��{dD��z�N$7��<���ۡ�)�����/�Ʈ��b��a����;���:ߒ�VzY�f�*|b;Zho�p)\v�n2��V��IR�i��1��}�,f��*�7�I�;ۓ�[@5��	���1WZ���C=0n��_�4�.��5��D��;g�ϳ�5)�H�duգ�)��L(z�)�@Z  z�Z� �x��CN6� 0W���R瀝^C���P���M��qz����z"�X)�ecy�n=�%�aZ]J�yG}+?fgF:�8�:H0}pKPwP�B�.G�̛�)��62?�G�f�w�\׎�!�[� ���M�����sA��ꥇ�k�+�`��iwMwl*o �s'	=Y� "�ƀ��7���|%�!Q�F��X��'�
��i�s��އǗ�l�7��q��%/�8���a,��"�@�)�x���'���$�B�|y�f��`t�
�%W4Vj����ҁpJ �::Z��#���A��{jc�P�g{^'�V@�@Z��Բ����Lq�����G�K�vK$�PH w�:Z}���Xr�I�nɵF���Ą���]�V���'U1_6�����f8̥m�'	�� z�讖�$��eR�Q�A�4��{�����X�p*< ��s�%�q��T�d!����	�{���v��K����LOX���R�'�g94BN��j ȃ���]�*Qu�D��Y�)ª�0:slE�Oi#�^�^h uq�<3ֲ��Nu,�L��CL� �Ta 7S��c%����g2 ��
ԏ8mKq�k�ّ�N)1��\���I_���ʲ��N��J"�{�q_�v6�5�z�A��hM���ww$��骑�S�Y�v7�����)�}�o�J�4�������̒�����L��?�5�hX�;�n�8�l�x�|aq{D����$	y��v�ܿM���Ԉ��5� T{�i�-�-��p�t�Mmӊ���8f?AO2+���ZKS���V�"�{a���E� j��l��Ó̧�BݘhN��=dDGi������1ǎ���kͥE���Sq��È[׃�d<6�[J��Z�k��0�>x����A}P��������\S	������V2��c�2�@j�_?r7��P�����|��dP�W���9�yWgDJ�3!:��
4x_X��}N^�pox�?T⼳��K�T�h�=P��҈�cpE]b^v��U ً;����r�D����i��U�qEd��;�������M',d�����ɟ������R���$N&�>�ױ��>�?���
�+�bD��f'�a�.ٿE\���R�̈�@r��+��9.s�������/;��{$0�Z�v��R���3C����U�|����_V�� Jhg7�P�Λ�7m��b"vxڀD�t��Qg���'tp!�&��J�ߏ�!3	�՞�5���wW�(M@c���g�=+*Ғ���_Vݪ�L(����z���z�j{A���˸�M��;�k���蹬@#s�w���}Y�i.CQ���䔚]	�2�\I檠Cl ����?��ȭp��rhUǇ�{��ء��-��"%�yQ��d�)<�t�齉���oO�#�]ճyc�/ʠf���c��F�(��t��w�&ɭWl�
��%T-��C8C�j�����ϓ�|�$����_���Xa㖷�po!�{�_�q|�M�I��(�iF�٦�1e&Q�g���Hx~�����B?���*kO�Be��i�j���z������I>/��:�=��~��������TO�3Bt�����D�N{�rFD]a���rk�^·����kHͮ���~-����ȁ���!OCT*ج/���ڒʑ�R���fd�ҫx���ʋ4��n6�0�����T��K���c���EOR� /�f�&2e�� �F����j[X��P%E���yf�V�n�`��Yb츫�&;K���"N�L��j]�����r0�4Qɤ�>�\y��D�p}��-L�e7���\c:��#�]����{.�^S5XE&%�T�U ��(N]�%k2�L���É��ߐ�:��E�4�J��܍c�_�{'E�`��S1se�$"����	�A��lz��a�n���hÓbn�|�)�m8ޙ�@��A�QT�CT����n��c:7q�Ѳ�����j��I���Fo������a�T��.���Q��407f�ξ�����1E�d�,�*Jl�ˁ��TV�-��
�X�]�\n"�~��� ��;7\���F[��9	�X��u�:���0:Ԩ�L7wfb�ԟ�*A���#{���|�r�b�ܐ���'�G[�T��8�N�����4��q��Bl1��\�i9���EĒ��V���6'nDp�Ir�x�Y�߷�3A����������)iY�5RW�����fr�9��=�Ƙ o�%B�ok�o�#�B�4�3��f�\^rpB5��f}s1��n�� c��Ԁ�N�ayʡ�0���٪6����x9T�|@�Lċ�#$o�Fs�Ȼ>G�h���93��I��pu�����+�w|`661��� .0�)�d����G�8<�񟑏ҬC�����W�洼&k=��߬)�ư�x*�E7�'Z���!����K��5�[Bs���v��r�������3H]�܉��Kt�AjIƀ2h��1�Fā��+�IҊ��Ak0�d���F"n[v��CY���8���~�J���f�\���8'������+@�j�b��"BW�-i����К���V��w����i�i����)�:*N�V=�V�\���ՊG_N���w踳�?�\}���e�R4N�{�[���N�o��>�,X���H���pD%3AQ�)���������u�����0k�`�]�z�;Z��{U���RN�T�ĝ��>���	���=�[�?�I�BD+�R���Ŏ�C��\���^����D�%���.��'jYҐ�ʩ[e:�.��~ܔ�>t�Z�ɺ~
�i$8	��e�GTT�,�Ԓ`ye��Ĝ�cQ��� л�T�6��q�Qm�v7eppզ�|�DwN>�Y�+OA;O�;d?�����z�n}=�&r��K��	�H)�m���`q�|��l��>ݮ��'d�~z橅����#���z�̈́8RG���b����泌�R;���aq��C$�%��V;�<	6��z���B����@�|/Q�@�4|g'��;$*�zdz�B�@�mGA�e顳�Ϳg��������Q��zG��?�=g��N�c�idR�Oo7��x16\��,H��${K�# 1�� HN{B�M����K�2o�.V�Z�o�K����LM�im�����_Tz���M�����3��^3��6�[s+�/t^ �ۭՑ�L���L�W��q�  M6�}[tGƇH��֑>$�������|N���y��)I��Zd�n_�/��f-0K�,�W"Y�>�H�Qj�V���������u��fa<�����t�/�ĸߚN7N����s/��9�쇆��f#��OXR�M����(�|�_��X�
Nc!{�\
ō@x�NM$�Ṹd2R�����@�m�6��z ����X�?`S'�3Ë�]&��N���f��C�A)#��&�)E�w{�Ll�)��Df�FLV���N��V3��@1�ǻ��؝�8��|f�8,5�����ҭ�J���4��> �s�G�so��
<6�r�#0��$�F�H��˺+� �Xؤ��$ܨ�8$�'��>�����u��K��j-�R���ҎE��O ��}
;*.{�U��=p�ف���[���)����f Z�u��v���/4v��Tt�R�9���K']��(/L8JI����! &ذ�l`��������9Q����W�g�8����ĵ�<�s�rF<@G8|�)�o�N���,\8���SU�H��u3g��}��E� t�啩H_��.�Ȩ\≀��B�_G)ED�/{2�0{��P�I�N��Q�o炍�
+vd7cK����&S�4&b<z�$��i,l������`��TT�n ]�F��|zx���y������A�M�=����5�����iI̾�7nƲ ��G����J^�%��:�H+B �+�ޡ��O�u��܏]~����G%2be�JJ����t�{�`̄�,����ڟ� Al�z��+y®�H����ID����o6=F+�r
(\)��JP#�.f�r�!�Zj]d%+^�p�h�>8 Im6�9Zk^�oK�l��TP�Vn�1,��'W42��Ųq�,�_,�1�������=y	�; �'q<�Xho���ڌ����}Wz���A_��K���⊉rF�~�w�1ږ`-Yg�5��u�!�?V�Zi��~�J=%�3�/<�$�i���
j�����󴉉p�Ҧ1�n�̙�4D� �������h6��z��]�H�>y�n�O��T�ٺ��$g|�`���߇���}�U=/��77�<�Ħ��۳H�\�Gd�dʕ��>k��B��扛# ��u���i�T�$�a9[�7*T�EH���݂�&KC9��&�?�s�۸���|���VDc�v�ҟ��RU?I�������q|A���>�=8^�5w
�D0o�ـ��D3���z�e�ib-A� ���7���O��@[��R���}e1�r��f
:%��P����N2D�a�)��Z{ܷ(}F�EO�=�M	�񅉾x�3ϋmc������5�l-�� o':tql��$�Mĥ���߭���g2��7Ç�«`�vҟ#���?�s��1	D��`��ߜ��]�X9ol����X��"����9k~��\��1�6�D�;��9�	>R��Q%���Q�m�@���?��/����m�Koz�f� ��V�u&��$�S��*o��	A<�Be��R�?�Q_{KB1j�؈��$JW���9�y�5`>� w��/��x���¡��������,�s���0X�W4ҍ���R�Ūv�ҹ<�pd��ȬdY�w���wH���4(��D&����l���Y��8@#\_H�5@foa��}�q���� ��o�׽����A�y
$3�3'��%#�.fg���ϣ��pѤ8�h�REP���G�}�kK���u���"��@�V�y�9<B�4�J�b��e~IZ)A��P\L��QC�]�̞�L�% �0����o�Lq#Z_�n>3J�)HN*H��O8^g�ګ���6��"�0���}�tV��{������UԠw���o�4A�4if
X�-L�bq�Gڑ	�ב��}�X���(����7�H��Q�!>%!	���~O{�"5l�A2�h|��<z�T��6����K&AI"^�e�F�Ļ��I�l��J�d6�i8.Q��]�DN[a$��1����Uo?I8|�̬��Ҁ����ԇ��_#[�DI��*��0�q�-秌#�Κ�{^ң?M@h�P2�8
kőRH0�4c����Iʈ����4�s+
X�o�H����̨�~˖)f�o�G@�H�m�f�\f��M�?ȹ{�w�b��{�)3.�h�]��V�p�������6Z��c�ת��}sE(�;srH��e�!�C�\U���7׫a�� ����#�ӓ|���ô�o̎�p� �\�?�
:�!�x��y{�XW��keo����Z�J�L&"Q�l(��58�$v(�,�۞95M����� b��d��5)��d�ÀP�)pf|���λFӭ��D+0֪���?��<�p��.�R��Sqw���W,B�4�-s	������6�9E�Ԫ27;�G��c$��+-5����\����:�bu�F���e�.\�����y����l{��~��Fj���0>�Si� �h����
QǙO/C��}���Q�Kc0ַ�="՛3�=���6�rø�ˌ������t�E����h3}NE�!#F��;P� �ei�������j���9�]E��aL	�i�N-�FXGOx��2�1��=X��zt��}��Iψ��K���L�x`f!=n��v�~؝�[���"c�d�$�|r��̼#J�ޟ44x�i�!�]j�(�+؈�*� ����;o�a�?}�X[�ۉ�-|��N�nc�;M�����b�i�ڏ�k$Ȼ��!�K� �x� �����IÕA��%��e�7�����L�@�L�_˾^�O�]e�B��f�L��.���D�n24m�������ǂ�Y<��BB)*?ci%\���{X�_�@g:8D6�}��f�Q8��?n��*����1c4 �����5����M�<�CY�]yr�G�N��fS�iM��CCM�$gNٕ�X24YB��=�[s�Iߝ��A�酛��r=Y4�/�i�V6��[G]#\hٳ��u� +����J8aљF-��w�����/�C��y�y�/̞)�J��Z��V���jل<��8��Ȇ�Uq�\��P��DD��o�v�R;�y�D����`��D�cH��8�M{u��F�U��"����_�[��%<������zRvy(�N�Z�v�A�?�&)\Fǿ��Y�}Yi����v��.cB���M�{!f~�ۂ�kwu����So��6��ݴ��7���O�
�+��ͮ|��}�jإ��]��Z�"�0bt#EB�
�Ǥ#C��v-�P�u�k�]��'�P����b��N~�Wۗ����F������p^/z���,��� ]������s�@Tf>���~������p�d��+�ћ��(�T�P�U���U����D����b�4G������uCb���E�RB�fa60�6��U"�%������%�r����r��k��\�pw�x*Å�z脅e-�=/ꀽW*� ��r�0kqxK���/���[��q��Q	��{�	�Ć��et�v)M�9��
��.Rfӎ@w��븗��Ă�:�tT�IV&�(dXFi�)#�R�7�m5q��[�'���9�O��JڤY�i��.��Ϸ�=��O�Y�������7�'+�+�Zߊ�[�C�np�<\)��@|�z(|��������Sxð؍���OdZ�.5���Sf��?��P.^K�X\�pF� >�Z�ԭ�oL���T]x�k�G�x2�.w%M),���2 �ۢ����,ZϽ8�b-�g��-J(��VOǟ���~Oaؗ�0�6��2;;�g}��^�@O��	��"b�k@�1��|����R�B��k��z'��r������5Nk+r�[�Eἶ�p_���{&���zt�>�h�P�2�#�����H���!���Q'� ���!�O��1i֫|T�w��!���z���dz(�U++�p�	�OV](�B���w,}"�4�|��ͯ�e�Vנ�h��C��QY;�AG�p���G
��!m���*yE!�V�1��Eں��ɶƲZ�ꮕ:O�)���%�K�A	�:�=�L��%g�B!.d�P������BD��w�Q��`b#��׷�'t^�.�Wd0��i�Q��)���"����icǷ7��D�o�Z���]�t��/��Ϲ�;��Ao=Uqi�m\]����K1��}��t���A�z���Y\3�U,Xn'�`TW:�G�ϗ��\�)��on�銅»lm������p�4Պ�މTY+�FMf��Pú'� ֞����Q���oOV��K�f�#kg�����J�vF�3@ ؼn�Nt\�*a�ϵ�dV�?b�5�gȜ?8��f*��[/`8X�(P��3+yu���`�C���:�Vnl<��|�3jI���j:##��>	��Fƴ2�<��e��.�2������#��W/p�����bA��i�T\ꊽ�o(]��t{��*�x▱Qj5�"Yf��O.��ڴ62TNN�w�/��a+Y���(F�ݳG�H�M�ڱ뮢*�D�����]�������E�k܂���1⧮�a��r��4a�^}�ij�B�x�}@����D�"n��j{q��Y�R�VA����j1�h8%ײd={���r�������B<~�l�_�kj|��Za����9�,"��C{ҕa{�y��2pA��i2��i=7�uE����m��,�A�9���Tt*��L�a�3uyo��a<B���J3Q��#G��72��,��b���p�]y�G��E}� F���Ĺ��A�EA�؟���뭎s8�Xw�k��Xv�FO��{�>�>��GC�����	�}����*k�BL�ֺ�SJ��7\Y�/W��BFd��A̡�`�y1�3��ElV����L�Ζ�����昩�LV���z�Y����h����7i�+����Z��UC.I�R�v�����B��%?V9rI�t �cZ#����>/����Rr�\H�l2��_mn�'o*[UY9��I���:*�C��A�[�r#��dvD6�B�B!�}^�C���Iqy���� vr�ն�]ʷtoY�Y/�3+Q�ഷj�}j�<oPӏ����5CSc�*F�j�TԚ�����JY���͵���>'���y�X���U�	;���]S1�\՜bil�� 3(�����p�����-6{K���n�#5�d���v�r�T���G(��a�2��d1{L[$9C�Y{��I��B`��?[!w+tr�l��y^�%�,9(*z��=�B%KH�<�%�C�؀�&s:�����h����3���˂�Z��Xf�k�ˏ(���A(�+pq���Y��T��}��'iƓ��$+��Aw��)<��oh�fK���2�}�]FٯAgޤ�#qik��o%dJ�X������]����_�V��:"��%�k9l&��H�����R��n��]L�v��2�{�2 X����P�$��kB8���Q;�C�`f�|Q0���G�e��3�\����N�B�(w��w':J!�ݾ�WIر*@� (���sDL3�p�)'c@F��7Yy����ة�g�@}��$�p���h��'�::[�ڔ4UĿ�X�f�7+�o�z|m�J�hq��l""���U���E�%7���H��롒�ɻ�e,�<�L���U�Jğo��y���� `܊*����wey2���m�Հ2�ղ��/2�V��me��CE�Ҷ�&}TU��J�^e�$�XU�ְ&a�a�f��ۥ�ܘ�����'��b+�92u���I2�}�w�!��,�t9��'o~���x@0�ٚqm�<b,�]���{���������TSң�(�%0 ����ay$5(�|�o�	�a�M�@����[���E���Hb�1��	F/�?�ƭ��o;.��К�~�"\��6<�D��q�Kn�J� =&�	�S���@(�t(]cp�N��j#h����Pp�oՅ�ϕF^{.-n�mP������#�����>��]����i�ޝ�8p?負+�q����������'v��i;�8����l?�E(����Y�pJ��h��v�ﬠ�+tGՃ+/5�)ԕ�MQ+���ط��b���,�$�[�p!���0���l�^*돜G��ƚ�lz!=O����[�ɨu�}Z�9��k��}ب���Ӌ� ��T���
.�o�rh�uU������2s���xJ�/��W����ZF1ؙ��{���=�Wi�(gH��2���|�J�P�W� �rXJt/�sz�A(���j����;oM���&|m�1�����}'Q �0�Y΀Tyh$��o�@0F0�˷Tr
�ւ�/fy����Uo��R&��1+�VNTBWՃ�{Dj�w��fR����ˏ�]�@�c��G���~�(����*�����%4�і��ǒ���P�;��Ϫ�S"�������F^T��쾿�d�j.���d���3U� �
���l�}Pa�B����歴�I�#nP>J>//7N��Y���Om�%*h�
�;uX���"�V��&=��1�!�oQ��)�u�����C�,��,�v�/m/Ԭ������]����؅?IV�'s+�D��`�vږ�YU�}�=30��Ǹ�ʿ3s����l�����:O��Qaa����\&�Njh�r!C[(��*%���R:�%<�w`͐P0FT)��'Y��>�`�O���Eq%+� /d�x�����;���ufk53Heҭq���W�<�C��W��B:�-2�zR^�Q�j�?����5���D�zȟ%yyx��S�֬ڸ,���yM����~����Uq�E�E8���eh�}�ɾ�C2s��|��o����z������D��&Ԯ>S�}��0�e0+�=�h�bQBa��f�L	�y���L����\��\ul��=��m�nD��{����ȦM�F�4O$g�DPs�n�h���4��-�q@�i ��E	��t�m��c�x�����F8��:2��8��g4P��4ߦ�U�˨\P{	�	�'��@͟��z{IYS֨jZ;�e�a5Ӗ�4�V� �v_u6����+��Kt�ck�� ���z��]`<��؟��H.�O��R)V�'��Q፽�a�qe1�$b����9Z��f<'C�s`�.���*�cA��$V��T��~��˴�y�>ۇ���r�D[P�mϫO��e��Aa�f, D���vl)Iی�3=�� ���
s��y3����趝������\i6c$���x��L�NY�琮T.9� !�^q ��A�"O,ܵ�N�JC��#�7E��&�� ��$��3$ύG���$@�?ǆtV�K�H/I��Qf�:����N�K.J`���KH�D���q=H�^�x)��i(݋QR�rT��ב`��v\`�@�Q��+�(���
<�׈���:�.�h��t��#ּ����@rq{� 0d��89�Q���[�q����$xO54��E�:�Z�[��-I�Ku]W���L�lO�ms"Dn.|���*��Ie�GR[���'TkJ��0Ä)ܾu[��,6����]�$�,tU>��*�)�u����Qd����^�SH�^S��p@({V�^����� G�E|����c�����a\�64�k���cM-D>�|�L0�pp������Cyڭ�/�æ�VC2� ��B�K��.�Q���xΑ�_�]��zg����J!�Ѣ����Mډ04(h�ۈ�d�CoM��x��Zk�(~���@�#��5���ᄟ�)L8�ȱ���Z�=�'����e�ϢG*V'm�RtT���&"N���8�L���[��Vz���z��$}}�]�/�p��f���|��(׳��2$_%���A�����&�y]��٠KЅ�Ixi̫��k��'.FׁIC�����"��d1I���\WegV�,��*)蜕>�<�������J���y���-��4�gTS�+���?�E^[FD�����)�ژ�j��KU͠~I��؃�\I�c2P�(�U�S`.#a��7!��77����^׮�߻Y�Uc�/��ֈ���.��Py7����ll<�&W/U6��������;�H��f��a�E>�hbT���q�!]gY���.�0��,.�ܟ�\��E��,��v�z�}_����iC}"���)|�dbm��Fp(���I���(���B2�>�������N�q��ߩx��3�������P�B�����{�v^~�e�so�԰�{!�,s�)Q�a%_�G)@[}�S�����t�q��2��GX|��o��s�&�Y_I�������%��d>��?��ϪV�p�r�G&V-ᮋ���S��гp&m�`5W�$�
F=`5l<~"�\��쨍�j6������*B�e�}(�����X��[w"�p/^w��{�הTjz^��TF��)�dr�:�
��d��#�Ԏ��B���pB,��]�uv����0\3�0�XN�1�n�.�1�L^�Y��W�浺ǂ��R�r��_Q�40���9�v��s�'G�¤G�����8(L0�66o�yk,�F��(��s�~?v��$\��`}�37��L�����EB��z���eq�j�"<�q�T�LVX��:�ˏ����0HX��r�R�%J�q誄}x�qSJ&�|�0�}a�I�L1h/P�r""j�B0�;2*/T8��4��N��l���Z%¹�} �]��^����]ˆ���^�,���Z�D�
�-בsW��r:tv8oJ�2J�]꜈��ߒ�V5����[4Q-��`F�<�:ήT��J��xVr��m�,�n�H�Z6�S�T'�Z��s�	�?[��c޾p�z瘵�� �����y��f�6�E�߅^��{-+?iZ��1���:��+#�1k�"��*Pu���rED���D}��YE������tB�GcbtTD��{�i��m�+ڻZ���_�p��}�Sn���w�^c��b	j��A������z�.�d���Jw��ҭ]�^7��{Szs�Y�P,I?~&3�� �C�C�_�����a�wX�<�>)�d�~;ɞsh�K�p���ծ�?&Ǻ�Ҍ����b�Bp��� j ��`n�����.���|,�JwFu��m6���s��wsj?�_&BAez�B�yeLW/������g���(���ɸ�f�a<
F���ʊ>�KZp �Uܳ�-�����r���#��[O�T9�KicxnzW�]�ow�}��Q����<�@��v����o�Q�� �	QP������mM;����c(1w��Ĵw�0�Y��!<�L�3�Ʉ�(�`�U�����-2TO�I�nw>���p��������8i@�w�c j$e�:Vx��bѸ��iX��*��q��/���	F������׬=x�������+lm�=C�u�N��Wۢ�ʖl��0����w��n�x��b1��{���%�Q����t)�b�q{����[R�fV�;(��ˢ�:�/(�H �3T�FD4N�N�~B{����<��r��i�����R��}	&a+tASSO��A`CN�O��F�B��(�üApE��2H)���fs3�,3��'����ƫ���Ehy�Cr�r(��3a1oI<'��~H���)`
\HlU��"�2�hؗh�h ȏ�]�X�V"ؚ�E�F�(:��w2�%%+ْQ�{��tk�G� �>B悝{Q	#�)M�0�Ӳ�^Y5�l/������p�xv#Pݤ�M������� @wt0����c�X��J���F��j���=&C���ߡ���p�w<d#ڈ���$R���j�+�A͕��AB�����m�Ka`<���5�
�$G��Ĩ(��ў>Z��?�?������.��7�z*�C�r�˚~b��������?�\J�|w����`0OzH���I��u�)��5��׉��v	�vE�89BXv�
Xa�o*6JMOƳ��[J66����׽M��$F?�ΈI_n�/��54��C�xA���~ 45�'vii�(K$��h"��)Na�>�"��#M�'�-��D���W�2��S�˘�w�u"|�ޙS>f�L��b�C���/�^�d��O*�m�P��5���J��v �p�' \L4zTJ�|{wG敝�SVg�m���m��T�E�-������Z~��ͭ���������E�z���_"F��4e�֔��H��Y��,!\��m���:�И��Pc��MèI1Mά�	ٷ�m�2k�%�%1y�q-�����˩��G��'Q8����9�L1z:��B�=eOެ��Z]�s)�hW�kg{��b����Y�r> ���}�5ΊW�|~�E\y6���l;7��Q�Y��Y��F3+ټ-�åEO*��!�B���?���p)UZ��V��~Ki�~=4Q^�s�e:��8w���J+5Ae�nz�E~8���cWz��v�4�	�n��F��]�6v���OBj?�:)@4I�z#��&H���!�1N `y���dZ�J���k�8T��b6�#'|�
��RP��Q�<?���J+�*غ�|O�bXK�?gZ�����`D�s���?�2��^6�_�#��R��nF!���JЀ�&;%}�^ӏҝ	.K�1�i2��j 78ʄ#a�H䫎�*����9و�06���O���%�+�Ld�G��i!/U)v��j�?��cX�n���ܩ	-?�&� ���ғ]kV� ?u��iH�N	��O,�Me�Xt�C���x�^��+�~v窊8�*��w\��(/#f>�$���=�/����3<g��`Ѧ�ӳ0��z����ԀC�J
��ȝ�p��oG��u��Dvt��N�-M�s�T�岞�y�y,����u�7]f��uO��j~�?W��¼bݩ��'õ��q�,X��~���!w"�C\O:�X�X�}��+Óf�ʀ1�h�{�;�6a�d�k����}�����'�v����.o	J����+�r������ȋ���&���󼁙OW����D�kM>��41l��Q�wBz�--������ڡ*솼t)zH�gah�<l��+���×b����$�߫y�5�]-��-ð�cү��c�*z�C<�"Y�C,�?0 k�vn>��mP`�5/P�{��U�����7�W��!V'�+N~/������;���I�1"rR�x��-@���-��;
�O�ܱ}�4�F!;5���~Ǣ����X�L/�#)��i Aqj.3��B�vx1���9�m����@�U|�@�ӛ�:��_[�s�#�`���u �M<�]��XK�=�SeԔʷ�\���$3�h#�vD����_՘�Y��\�l���!�Pmͫ8)UE����
�
,� �=�LɷT�'���m�y)V�S��u"r��n��ą*z��(��o;̈́��CC������Ә��]�=��ƲD������Y�}�,n�;�;l�MǞl��zJ۔���H��}Ţ�F�}!��/6�H��x�Q��~fp�����nj�{�u�l�\�LC���"��PƬ��Á~F]b��<��r�U7��.�p��z	],9��$�~���4�;�zPh��mF$���1,Q�Uݟv����'8`����	��O�#ǝ3�4�x�K%�{�G!B�y۾�j����W\�F��i/��,E8�/ߒ��1'G~�J�8��#'��0r�<�u�@����BE=��),���*�;Ӈ'�_��/N�p�����U0���mzOJ��AX�j� ���kDCM�+�
W桘����qc|�b���(�B��4�^��ܡF����(����U	k�6�V>�Y�+9�4���q��nbJ��<Yr� =��uc�7��SR���Z�}Oj'L�S�S�gR�7PI�o4{���ӟK�+�+�.v��se�ZR�f�=V��n9g��%�{J�B�EM��}������sg~��r!��D�!��&��|�$�nz�N6 P6R8�{�����1,E�D|��,nܵW��@��� �Q�jvM�Dy��zsuݽY2�x��?�w�z�og{,�v�[�i���l3��]�aZ��w���m�q�U�X]؃PS�QS9�;8�Q^��An*)���-��oZ6µ��nr$L�2_��v�#�a9�@�at�noanM�����|�W><����U�:?���óR�!�6��R{��s�\��Lf�mM2�ԩ�1���05�� U�Z	a�2�%�Q�b��e��ŵ[�����E�N3�%fn�d`�	�e4�c�ma�~�g�-�D�?��6��H��S'�<(���ELo8�+�,�i����#c��	3�*Gz�/�^�#�0�+�R9�=�H�m)^�ȑ�u(ݚ�am'�?O�kws!�{we
ה�V�K x�6�C���S������=��}�ξ�hf$���)���J8	� ��"�i�(�@�j�۴s�R�Kk��B1��M����5Y`P�l�25����p�ϡ�_j�>e��IX�3�{K�?��ok����r�7]�U���=Z��q��9aGhn�{�U��E/Ǥc�x8F�h�3�t+ǬZ��Xy6YD��<OG��"�e�x�B�F]�?/�3�wҢ��W�x�(���'��ď�	sE>���p��Ul�PB����W��?����W�&�1Lb�rdd-;v	��\H�;�p7�My�t6ΜS�>tç4������kRa��Z=\�	ca����O�z����"¸h]R�p��^��Q�#-)�l��n��<�ݢVZVm MK�'`cU(�ȥ���E�c
���*`-�݆�8G.2�U�6��~ ����琔ܣ�����m(�AL�'� ��M��7
|�l4�E�*c �C���l�3+B�7@w����r�@09ܬ@�%&a��W��^���h�]*.O��4�%a	\�n9!ktXp��dKa�U2'�����<��o-̕� ���λ�[���ڀ�}>D����cN�b+wȥ��.�;�����$�����;�)Q���������a]����>��"n��~��N���"%7�g�8��3�6�N���⅟�5{���ob�n%��;씯gbS����9��&n�EioE�-��؛CZ�7H̅wgR�)fA� ;�����-�YE�ד�'��MO��?�sɳs�fg��$�z����A���q+s���ЁL���&����D���V�K��'����u0�q
@ie�%Ü
F�_*hc<>	Co��u�n�x,��>��W���V�'�D��#<tu,��<���Ja�{�'�[Z�/|Ɗ9�8��5" �d�!�5�Vs�V�vb�b����1´������h�e�u?�����=p��첃�nl���X�> ��- gUd,~K�y��桝�U[�w"Z^c��Ǝ-���
�wƹ���#v����=�C��fI'�3�,#���EV�br ��on���5��m���ΰ��,�O[Y ��,˹9�}=nv�]H8�C��2��-�7�f�����om��Ol�������\14���.�^�L���v�ĸ�������U>p�Y<�|����03�Q9:�X����f�?��o�'w�;����H�zB�y�xV�,4՜��T�/���������d�.{lGhr�������8w�~�L�O�Ԩ�$K�>ա�&�����1��:����/�XZpy=����6��_Yw1Q��(�VQ<����-�0S�h}$'�����%�&��9Z�UWv�K�ֳ}���lu8���}x<gJhc��@wƠ��8F�k�D�yѨel�:��[�L��>|!�FZ,��W��,	���j�F_;<�`ZR����$�e���~Ĭ��H�RI��,͐/+���eU	�-B�>Oj����@�e��=zZ"�	�{6d�o�#5X��Ѥi�\N�ЁjKAN����>��2���'�T�uͪ��8m�<�#�����O��[�����7�)8����u"��a�KtT�I��q�<�Iem�[G����������Ie�C+'��/���M��	$N���L�}6hMF��O�zBx�XN��GO>��]���X����g�6�ۍ�p�Ө-���Å�2�ec�O^s*�#����u$��,�H�M}ӹ-�F��6�PH&H����M�U�㒴�alR�'s=��P3�.��p�=n��œ�T���S|�m�j�R~˓�,��%�-��R�x�-/�8T*��J:�V�l��!�if+�X�?�2��6��he2�k�j��H��PN��$��34�9IЭ?��̖���Ǌ�b�:�C՗�˟��������ߟg�IX9V�,}}
��W�7�h����|�4��]p�"dǎ�BY)�n�O�#�G}��S�V���򧏁��,���;��"�5�?��*2#w�Pg ���)Cjc
¬�9�P
��t�����]S�5�I����B���؀_�؃+��ot��.'�Ό�O�����P\�S�hF �nEPF�Z���S��bE� �1w9)C#��G����zL���V�4Uy�8��
6�������r��Nz�A�\�;��
]B���ţ����ńE�Q��uZ��$UP�'�ahۖ/�_x������M��j�y��B�����5�a���ڷhh��,��fg4hܸ<bH�����qw&�pf�<�!J	�h=o��vk�P���K�
��w"��N���Ė+C/Lu,`�0�����}�[_��c�'-�	�R����OY(�ʁ�a#�ù�u�V��1�b\+ɵ!4OT�����BL�ՈQ�N���z=i~u��=�S)�t增�;r�\��'y���l�v�U .91�~���Y&�)�Ț��#z�%J�����ֹ���[�����}�,���t�z!�{�
;�����W�۩	H-��n�&����UtN[�j���`�
i��� ��9�
�~�"l_�46TΜ4�	�	
0��@Ks���LLU�H9i�D�����Wޑ+�U��J��}Z_O��� ���m;��<r�Xd�����cp�n���[P��(s�3-��2Pz�x�8O��=:�n$��OO�f��=��7���+��n� \�_Ə*�E�*����מ~M���\䕯X�d�Ҕl �?��Q�Jm��ppOy� �~��Ȓe� Kx��TFw�� ~��W����j�4s�ޱj7}+�s8�ږu@?�C_���~�!N�aHp=��b]��l�6^i���R�w��d竗�A���_Z4���B.��
�Q��� a \':�2��<���x���vdW�꓈H�z��`����F俓����ӣ;F}p|��
��3�5�
��2g���^��"#����29NK�'��H� v��n"���wbU�v�q�q2��-�O����=u �:%�ԧ\K��Ȕ�ʼʁ��9��`�H���c�d"d"�Oc�K$��`��}�J%Z�H�?*b}Yj����J�!U+su?�h�z,V��\Œ�0���w8�z9�O%/�>!�|�R��:=���p�&#?����t�Q���7mD���m�Yv\�Ph�1��FMv�c�k�ڛ�=�)É%���Ыɶ�)�[�]������rxy�7�t�8q�Ǫ""�B^`�0M�~nakɶ�_���N*�P>��J4跓\&�k g>b����7+�Tn�&X����m�Tl���bI��og�3���t�ۗ��k�P.[��$�8�%AZR��~�i7[���n���s�N�sO��Ň���S��I
����=���	E$�w)�&�p��?�粻����"�����Cj�[���Iy;؊����<mc��+{��b d��}�![�w;yJ��;�@��߻�����˅��ݩM�����&-�.�E��G��o�ĿZ,���_�Q{���<z�����l�b5�M��-�jgk��i��#x�e�҅P	j�]�v��t��Ti��=o�R�_����?Ǵr���ӌ�7I��_C�F��M󚉝s`�K7�H[h�����&� �F�>�0��'�yG_��AWm��O����66Ziͅ
L[�ukgXL%���`/WԽ���x�N�,^��c�&�3��Uv�ANG*�#_��v��y2�Ƶ"�?oC��_�-)�����(f������1�>��ZV����i�L��-3�'�4� �[��a���P�5f�er����R�޼}.��
�<�48�r\��'�a�&�����r1�0U���U��_�j  :���*�x*uO��7,�t���Sv�3�MX����4/-f��&I��97���!բ���@$�
}�V�I�8���#�:l�v�(Rs�Z�/WBH�lx�"R���@4@l�$�*!u���ԟ��"+%t��{YW5+�]<�i�8�ɹ�Lj6�I�ؑ�O��m��m��G?��t�#I}�/��3Pm��-M)+?x_O��>�A`Ѣ�[YC������ ����<.P*\x�!�=9��9&<ýQO�q�Z�6�
u�V�A��|ZR�_% �o]:��]�l�6��%Q���	7[`��|f
?{}�`� [ɨk���S4����o�|~���������%�F�͠b�fj�O��BA��bϸ}����,��׊j��ivP�Fo!�r�D6��3`���F9��f4�J?w�i��t#m+�II�u���9��k�#�G�.���F��e�M|Ph��������w��
�x��
~�+�M�D܋� kӹ也P)�Rur� �Q��P�v�N��g�ˈ⡅vh�8����e:���5�U?06�|�%I�g�W󯪽<�z1=�&�UT�o���g@�qΙP	��"��@zW��WʪB�h�b�1)�:?�.�6:g���4�*�����s�y�g�I0�̗�ytrY�~ث0|vb�(��J�����n����n��`y�A��o�@&jD�n?�/p{��gj@��2nB��lj,��6?#�(h7ہ�%��E���u�k���^�H�ӵ�M)XC �Я�ڟ�L�=yWJ=@-!&�����5,B���Y�Z�_�_ 2��v�ǲ
�W��Y���6�r�}��D��E�H���7�-G����G��ߋ�W��M�U�@U�)��.:+7�&�+e$�b&�	��~������י��َ����>m��Yچ����xO�\SK��1w���*����
K�*�Zյ����p�Қ�՟J�[�y
�XJTS�~u��b��#��(o���a���b7�|O&߃�@��0�<�Ŵ�Z��3r(�2;ę�q]'�]|�*��+%��Bɐ��U��v!�����n��d��z�y�(e밉��/���*�z�~�ϡ���<�����ԉ�HI�Q����j�?�ɷ�p���6�:^]���v%��6�� *Y�TQg��:!�Β�T`{g�1�b�W9���@k�����Y&��T�}�|��eײ��Z�A&����U���*Dm�Bvz�(��R��T��Juk�o�Ğ��J�y��
�U~�TE��W�����jJ�^-�tPk�\��2��R��xI@C ��Pz( G�I�]�t����#;�1�+�@����7�~�l7��hJ"��U�Dx�D��|�"b��稨�,�Uv� ��(�<�ܻ[���{N��v�{ �u�?��z-�sg�Ar�/�(}i�Ȏ�{%z��]��V�P�D�����bx �>�$�ǘ�(�_����ߵ��{���|Dp�  Us<�]͡ª[
�#����=H��D���DF�1JZ]��z�1��X���R���$���i@�|�NЃ��C>������Pw�b�+���ǃ�v�'�ԣ��~�U"�J��cبA���YUN�F�l�P�	�0Qn��M��t�JL��p[U�桏����SF�5Y=k�G���M�ޅ9i���/J1��2Ɵ�+��ם�!IH�� ����^�7��H�U��"9$Ŵ׳X��ҥ-� 1�޲#������'�6h�|���|�0o����~�D@0 B�³bq=\���H�Χ�J���C\R�
����^�ԋ���=�s���	�o:�o�}��*�������?��;|�׷\������-8�,������W�����M`�������D����tǂ5.����͑&�6���� ���&íF� SJsb�35x%�Cԃ`䠐�L�y����q�_b�'Ir��=t�J�5��	�������ê�s��8�/��!x���W�+=�����N>�e�J�?����&����d�) (����\�F�x��6(�2�6�2�Բ�(iK��:#�֒RL�U��釬��67��B{.�kNRS��J�VtƼ�Y���_{��:P]�F�ː��ϡ��d� �SL#�a��[��Q1����7���&���A�z3�w�<º�������G���£=PH��sCQb��͒��a"�?�-�k�&u���^�D,�2�*�&m�:���`A�?U����n��,[��5Z��Ξ�(��h]$1$�n�3P]�o盬M�ݿt�F�. �A'��go��u�U�!2�M.M�=��`����5Zr\4qbw���ݱ�܄[6�2�B�^7�� }�3��#�@���{��1*c]^����	�oF�;���|���Pl����K'��Ru�lLd���{>��,��ij��AA�K�Zs�SŮ����PbI��o���ߝ��:Q(�7�<)^=���Z�a[�|/�6�ɟm�\�H���*N��lӢE�#OZ���NO�ա�ߺ�K`����T���2�S�A��n3�hY�6ح��$��L[�.��h p����
��0��D��(�SyE/�`�g�F
7hR� ��t��	�'a[���7'�L,I�C ��Ӭ��^��,��o�_��G�9�Ho�؍��½d�p�)�mO8Q�00�� qضaai��KL�Le5��Pw�[�f�	�g��9��'��K�bAǟ�k�H��1�j<�x�s+�y{��ܾ]O�t��U�2�%<xx��J �q� �d� 9(h.�T���[��$ʟ$qM��y˂�]�T�����t��ۚ���I�Im�&��B-4��@��A���r�)ߒ&ٌ���~y12/e���W���R�l�&���6����A\i����Ua4���'�eb N@׬6��p�w(q:Ka�4�d���pCC�[�u����M��<�SFRϧ),Ulo�Dzڊ�,^e��\��$��{jL�]U$�e��+ct��G'�_����v��8 ��*�.�@�1`�F�܎݄M*���\Ȝ^4����8ki��γ�d��M�����
!L�?c�!�̭ ���:W�@�����0i
�*0Z�O��t��ez3S�T+�Fy�Z����]K���\ߪ(�����:��S٦u�{w,���|�\��I���s-�4�i��/j3��\��'B����ÏO�թ����+�^�Ռ8���B�2e���ȑ�o�[�G��OѵI��ac^�k�筸qL/2�x����u�C��V�<����V���$����x�Bm��T��t�2�¡`�w�mk�E�� S��zƗ�}y�����٩���;#�2@��M��G�M��\����B�q󼙚1� ���3�8�m{X�� F 5yyԩ�n��X��H�o b�U�r[���Ǭ���ٱ������Ts���nD5��	�'C�Jg�J}DI�c�<T2,����^]1�w��ӻ���wLr�qD�f�W����Aq��{�Ęq��������<��X�5��~��[l���~R`g$�K�ᣐ���S�Ѿ������%|��E1�N���v�� 2h�ՙ���LR]����T�k�R^�T�{!]3��뇯l
�t������[#���C}�۬�F�e�I5�ط�ߖj��a�kq
���h4���l���_�$�TH��$���|B̨E8� �?~���=D.^쀇l����RNP�V��)q|�1��?}IKHx���b*��עT�-<������7��x�g��Ԁ)�S���֒�Y�p1 ?9>#j
����O� iG�A���{Z T@�;���#E����{��G���^��ܓ��hT-Q�XNB�sݴ��U�8@�a�d
�-��}��=�-�8�������Kӡa�u� �m
n�"�
[J~�9&�,��Ų�P��I��谗��Č�qL��*�+-�����׃	L���ܖ��>
4�[hsM4�-���Q�/{�L{r{}~+G�R�5���{_�8�{�x��C���[(AJ��u��-����tg����Q|�4�\�n�ř�¾�WoIJ��tg�G|�o�D ��O�m_�S��Æ�*+�������k��A�N�H��t|�)ɓ��0#|��`�eV��Ɯj���#(xO�V��L�����vROK�q!�#1zѴ��H��ˇ�쒓�A31��o�h���H
W�cE���0�	H�X�RZ��|�JE܁��Kaǌ+��U�(?�*�R�=N�%[��1�P������-jd�[�P�J�.�ր%_,��w���҆dv7e�}�<�Y����73�;��4�,KB:\B���C9	� d-d �e	�B��^�I,z�Y�@p0l��A�S�� �"x�}/��z}�u�S�h�TeBY���BB5��Tg�%�@�������R
�Z>3�����"!t�ܬ]	���>�$����@>"v � �F�4E/�`R�۽�h,JN�B��H����b|�!�Bo�A�%�Q���6�,��1R6\#�
�4��_i�!ו��/����$�:-�~��Kgt�5�!L��%ר^��/T�w��)��LXX?�V�#~^�*���:3ծ�_:1����Z墚�ö��L�~������G�{?ޗ͂=����k�Z�r6y2+�@m�<�Cy�A��� \6��15(��Z���%4&ৠJb#|��R�f(q;�)��M��?���o8Z������Y��rlX�(a�YERw)e��iS�i�#V��)�M�e<K�h6'���x.RL����ʹ	08/$n�{���+��Bt�E�B�2��,�Pֈ:�p��Yy�0�c	������fBu��([����=9P��5^��@Q�Z�膽��'ړ!�b�ʚ\�Շ��?��G��-�����M��E�t�Y���"s�k��ۜ�W�&6A�7���{�x���EA� W;t�����j
�G��ؘ�A �� �}t�/���0����z�g,ivJ"ވ����3U6D��R5�{^^wΠ~Y'S��;�ҫ��:����� &�0���} ei�j���9����j�Y�6�Ll�R�oWh�Ӵd!O��q]��q4�P��2Q{�JϽ��X�,�Dyf���򢁙���5���4�q"�I����+`��Y���<�Ҥ���������;���=������H��� q;�z�L���L7q�Y�'}���\{��ǅG[!�	�/�菩R+�8^��V��I@a������^i�բ�t���	Ƣ�����C��q����{-h�P���k��N���0(V%%X��J�:�k1�_Q�:�	,��D���F�5��g�gG_��3�:�&!�-R&�"{;��Y��
a]k�\U#�"� Eb-���!�~y ��&���F��}���#�*��p*K�7&�}zȻܒ/jNW�}��J�9�\`�>�W��u</�%�,�R��O�C�z{t|fҠLw�t�ęX��O��1�z�&˖݇R"���kޛg�w�:�Lo�0R �c�idaS�\?�R�S��T����w��98��㍾m�'���hͦ6��7���*~7�^�-5��(yC_}��U�V�]C��ϖ�e�)C��Ԣ7G�P��=��ʫ FK��p�s`P�jL+�R`m�uN�@	�ċ��Y<(߬mB���|��<%��]���<��7Ђ��F��<�x �=����j��P!��ryǘ��:?���%|��$�;�K��Y��T�l.�"P���l��q��F��T�G�48j��ѡ�v�OC]�i�&�t �1��H��Fr���՘Z"����q66M�Q^��{�	��>vZD 4�����NDܧ�wX�De[�d���S����c�ꠅn��2t";+K��� ��l,�_Q^J���U�X�j�y&V`q(��փB,��y��� ��ٙRs���
d+ւZ�jA[r|�����;�q�P�R�;��l��I��
w��t��.2��K�ɚʟ��� t� C�a�Ϛ{���:_O�4�|B��hU-H��{<�3��I9p8�ԟ�72:#���Lz(j"oj�e�x�<@>��33�+����m����`�6�GaQ���`Q�?��f�o��.W'Ǥ�J[��Z�	8� Nr�Ц�7��-���4d���LJ���.�ᚏñ���,�R��!�P��W�f��� ҹ�d�C���)c��ݿ��h%]`\��*M�8�����8=K�^�k��O���k�wd���s�_��Է��x�b0��*�GD����01�h�z�"	���c9���r6-O�z��z.�ނM�������V��������dX�H�^s�	gs�?�^J��@[e�tiS�3�1���Υ>�i �gE5}rV������*�9-J��G�}?.vi��pW�?��ɡ���7;�ӹ�
���ͅX�4J�������љ��|(�;>{�j�x�`95�����i=�rN-|���D,�&�|���H�_�8�x/����B觷N��J��qn1��$���R�M��>����� R����\�9�{%\�����9�Fx�2k��΄��N���K�	��kѧ���U���m���	`��d��,��*���8��T���w���-j�-�)X�,f��;���ު�����L��D�Ը�f�艹����s��G�7��.�F�SX��lN�#}/_�#�dg_��O�j��7"�~�o�C��˺$��>�,�T7P� Ȧ�	&�K��Zݬp������U�-mv#b�=�ݛ ���`{^]Ug��et�]��g�]�?s(���E�V�x�-�~q���h�[lQ���-��u�ף^m�zM����0�������hWK��t"0���߂c؛�Y��+��C�V���퇍WfWf����NSfW��w7�L�)ȡ9�s����mcȖ����*7��=Q&OƠS4A�T秈�Tv1_���Ԛ���U#z^ڕ9�.f�x�+A&�����L�$�n����~b"���͚�a���?��_�W���R�T�֤��)S �S�@�K�l&����3\ے��/UK!����L��.��u�%)��F��v�څ��
c�by��8�\Q[l�%\(��j4��E��XL��[��� 
��x�8��בp��"��U���?z����r���5;��Jޜ�"��*V�.��x��h�R��1,��'��^n��Ⓣ�^��a�p@��(l��#���X�',j���SZ�.�Q���{���l,?0?t	ށH����̒�꾋O�;��&���3h�{���Z��ճ¶Տ9�^z���w�i7�:O�v�CG��W��ƅ���{��s�qؠ��Nj7<�u� C�����-��h�Y�_�	�����	�_6���~�ӧ�jg�I:}�*ǵ����9s�@���YJ�J`�e�c-�6%�A�c�Y��p���%s��T��m���f����Cy��.繰{���Β�i���ն���^��:��^����-��J�rky�{���=O0�]���\��i�~��Y�p"7�'07������������j��<v�'����p�P���BĦ| ݕu�8�fYܐmW6�h�;�TU!�q�n
ɉ��=���h!�1�+�H<O�����,DjXS����A��GGWz���v�R5�P�X�Ώ��}�~U-�.�����[�.g���ycJ�{Y�;�T-e�{��`��l�v18^��ր�8����e�Ufv9���d6r	��zq�i3����zGꃣU_�o(��e�o ��(���%C��8-}�	��w���֒?�������DJ��J�E�-�Mo�� <|��Ιap)��>��=~x$я)���;�e�vF���/�L`�9hU����kĒ�G��1�?����o��Ӌ(�0j��������0���^p����I�G��HO�7{��n@u�D1,;�S�%/����T�ͮ�2����+�h)�-�s��23��ֶ�߈�ᓷ�˲���^#)� �ܥ��Nς�V��K����#��`���Zu�G��8t玟����@�߭�TB�劓��K��b���P���-l.EeQ$����`���ᵋ�m�a7�H�ڲ�ZPz�dI�Mr5���A6Ώ�ݝ	j�|K`�����:1�A3�k$���hm�2�����*V	�����}���4���р$.���f�Gԁ0s��V��i���S�CVQ�hZ����c��}~�����Eդ���;%���<n��(#7y��ba&�6P��7 �Nh}���]"=GN�}|k\+4���9��u�G��L��[歘%�4�If�H�D�/��~�k2��1���~&p(����:~-�5oI.�*i��$u���\½��4����ao�Ė�K���{�:�VV:��ۣj"�J#� 3}�Io��ï��b%� �2J��Ls��I���`D�FK2��!�t(}�AA��u6�X�]O�XҐG�G��"�}���gi!�I�T$��N��'�9�\��yx�k$-���0#�n2x�!W�z�|;�KFڣ�B�	����C�]Yͺ�i}=�8��q:w��`{~�/��e��*��3��Z�m��֍���%�I�RQcm�冶��nt���W?�.�ZuzɎ�����M1�@a��{��ǲ�����K��5)�5$�"��c��#t菬jߋ���Y='�����yg�P�r� k��6U9��7O���`�4���DH��DfړsH�_�9#��G�KAl�d������oI؁�jd$ي��U(u�`� [��1��b)p�� �����#+E�<^E�UmRj��;�ֈ���Rb�� ��7��Z!�;�p^��������r���P��2�gW�����l��M����bY��ۛȦ���#3��K!o5��ab�<pg����!��Y�t���QOjf6/g�wA�S��T�6c�7��B���1	�@�s��Lfu���хJ��9����w��S��.��%f�:�{�Ua�(W)a�iD�bj�`B������rX��I��
�ܨT�M�/BcB����l[x�u�,!v#'Oӫ"��^H5�5��+WRA�0�T����E�#�(���T��x�x�K���
�B�#j�V���it�(tK_��ܬ8o�j�/��إyA��`)_Y��^:���O����%�ڵ��(U:�������V�ܳ��	��?��sg�� ���-�I4;w"�"(CK0海��,X�n��/Ȝ!
��f"�K��ĩ�
u∔���ǁ�K�{�=U�TvW ]>:��A������]Ii�y�]s��3��n�	����r�k�4�#��Q@+.��B�I������to4��r��#���Fdy�0"?^25���|�ж�^��t4�u�B5ncV�4�����m[B�\��]����=p;]K���e�´�т�SKB�9��nܩ"��-��}$&aV|���q=�Ĭz\�I��u��[���J�J�]r��0y���?���Ӱo��4��_�A�Ti�Vc�EV]d,�����*?��Gr�:
O|����1���p(�gf�s��>O!��ֹ�����&�=6��n�yik�<m�-��p�\�
�T�(z]�DG�p�?��5j4ȍd�GH�ַ,_3iIv�R32��΅*��d��^�&Oy��,�S��.���ڽ̌ �����YS-G��X;)�-�$7v�ދP��r�Y�b�̶P'�5��n�c�7B�gܺW��_���ǝs[�؀ix5�}(fu��05Cx1z��E��N���g������>wo}��)zx�o>��uI�C��/���xŅ�^��,��>���^ν�e�s	p�O..;�n5ȫ<&��5����W�Z�^��f߹��t�(�X�e�Df�6AkGF}Ն�/O�M{L8�V� Ϳ�4m��;���ȫk�׆�o�"���R��92D��r�� :uA$r	U��~c�ڜ��>� �����d��Ȋ��Y��8/z q����K[q�
�l��-Y�'���
���4
z�<�A��B��㧟�d[���Qɥ*���ͱ⽔܊��9��������y�K�����a3i�K��O��k5�YjKY���ARݷ�$d��� V���������(�d���G�2��W<�r*�E_����P�|���@9�#*k"�m��"�����39���rq�zb)��S9L%�צ�Sɷ���e �i�2��p̘������M��)'�Mn���-aT���Z{�?�jF>�rzQ`*�[vհ$�D]K�F�.��~F�j��'M����)A ���O9���!/Q�;���P���I˔���`��Jp�B�i�n�~���^F�	����I���z����K{@��T�����hf,w���'��B���:!�N+�[��Ž?Y����	}���c��I�L�p(E�t��ꀲ�������ް��|�Ơ-@�}�C�#+�R1j��!������z��c��j�mDAj��p0�������`�_DI�7��k�9�&U���V~���q�������Z��ࢪ��}��q��Z� �Pyʹ�n��Eޡ<�
3��|�����
�4ق�EQ��p��"����Q@�[��a��`�]�l��/6)����.�7B�J��7�Q���K�'�Y�$ˊ�"%}�F0Q�Ѣ(*�d��*,{E�?칋l�N'��n�*s)(��$V��z]�E���G�ʗ�$W}�s,��&�Y��5�n�Qn	�,"L�<{�rGF^8�����Z~8���b�A���*[�H!�9���ܑ��Y�� �ٿ�$�|��rR��-._L�S%��8�O���qX��4�D�p���۞���;Y ���%]�����|ܒ��^fN3N��%��-��˽���!�m9/�|EO��@H��<F�[���M���)���_̲��E��W�ܤ~�C��f�w�����g���&�X�ع{9�f'�A���>Ҥ?*M0�%�r�fw4t��C<�U�m��uŧ3hB�f�(�n�g��5dW��s��!_H�T�C]p82r�='��JB*~N��I���?j���jlS���_~$� �X�~�G�`�y5qU���g���l�kA�0��i��L���M]����'��������Q��(
Yu9X�Cm�0$oZ*�2�L��.�x�����"��njm��d�!���\�Ve&�*<�N��[������<���>�ؓi=q|���vB� �c���AW8���|�|tHP���� |^�2��Q�u0�%]'���:t'�~Y6���Y��7���u<r-��o*ʍ=:ަʴ�zm7u��+[��5��}�g+� ֠X6�/��&�E�6�StX���f� ?@�,��[��^`d��	��{�,�5����Ͻ?#�}�����x*��ό=#^5���H�A�*"�~�'���IA a����:��@�'�3�y�u����o�d���+��a
0��k4�H�v$2
��]��uNi����7i]%�m۲�����6�������F��b�Ef�B >x����J�D��~g:F�ȏN�e��E�07NG�Os�����I�_����U]���ƥ�*�A�B1��q��}/�6��ghQP~���7v��� �;��W*kH���l,�5=�!�%8��vfXv�Ց'	�/vLF�:�ٶ��L�!�D3Ď;�bD�N7�V�!���W�P�5�CH�]q=�0g�\F��o� ^��`������xB�8g���b9����H���9&5�KN��<���?�AG
e�͞ޙvND���5�Jw�}c�D/|-i!��{��A�"��͗����Y4f`x��$���}{����
�@Nޑ��Q��ru�np�3�;�iC\SQ�.��Gkr;�4�"� �
�Ib��e({g�Ş?�7	�C���G��7���T��:�o�[�nX����W i9G��ҫ޵��Nݑ�D���u2R������CI�V��k��Q�P,CY/U�8
9�7E뛖�F*w�8���������D�j�r�cN���o�^�͹F�vq�e����G�-�~a؎u���d���~3[|C��S�����JGSOIMb|<�ۯ���	�~G��>���b�M�%�]���
�؞X��)�-Y��)�a��(2IPZ���f��-��?c#��&�ɯu��[j�gO��yV$j|��LY�H#�UU��� ,����֐Atr>�*H	V�2�Y����p\<-��^K��T���-j	�f�,�曨m4�S+_z��76�-�9�@���n�L��b����M||f����wV6�$4{�7�J��b*>[����ħ�I����%��K�bu�?���菥�%�`4����Z�r����S0{&��iK�?8TK=��ʼ'�GE#��{����b��܇���	ƹ���<�p�J�6:��w���'	��W�㷖P@J�YfbX] ��k�*�j<��c*|�H�)�:�
���J�&/�M��U��J� ,I�K�Ɓr�*;� ̪��$��'�$��eF��z�eg�d�
w~V^~�j�GV�yI�0����>���p��g�x��r��b�*��s��<��P���Wq/2�����Atl��%��sۛ��:�ޯIc&��y�D���$���|��9�/	u+�f�J���9��ϦPL4�u+ k�r�g���)�

)�S�<ǾkV��r6+4�6a�=��dR�S7С~����$@L��훋�T1�?B�I��q�a	>��`q�:��K���	G w�*�oX�	�Z�U(`8��#C�����1HGH�Q
�å=���]�q<�������ϛt!�A�6q��L�0Ƌ�r�J�3�G�h0����G1������ܥ�y�A��N� �A)�x�t�{�1!����Ŭ���"V ��^�ۭ�·�̶�����:�߰���{=���|L���g�~c��fb�}dz��T�G��r�=������=����9�I�)+�<@߳@�列��:
r��-I��N_۞���|u�]�Ǿ'�]��̵��üj�]�d2
N�.quu	?e���ӏ�����fM��!Lbyt�fl�b�4�BQ��o��țcУ`ŝ-�ޠ��F�E�'gSj��D�B��1�S�M^ybW��є�'�0��x�YX�T�\�ɣ���������sZw�v�x'�w;]_s�D�56�]L`�o�Rp�+C�-�t]�t�J^�ˊOG\���z�+^�1�r�Bp�9�XbHΒ���@*��&�Gk����}L��z勇!����D����ͮY�S��\lj��S3�Q�Y�����΁�$��y���C"!21��Ӹ$���,r�"��%���Hj�;z��Q��5��o,�o�W��
u����ľg7;F�9^9�ƽ0�.��*��vsk亵4�qC�����{'YWрf)�R�f�V��Е# �K�~���L�OV��r}CÀ����Յ�(��sUl�l�σhp�ĎSަ���3~����!M0��__D�~ႝW�?)�l�F��0�8�r�h��z�T�8���1+���X�d�[�2��\����Vӛ�d2R�E����eB+�F��������ǉ��2%+�<�'���e �GMC�`Pb;\��h���<H���@:�~d���--X�A��p&U����a�G����7W7���
c��/��*ɵ�4g�k��b�Rq�����	���*+yX��t��'�7?�QK��#P;�-y��+�H��O�4
 ��B{����
�sF���];��ۆ�p�7�s���d���vb���e�^8����$�?�Ե`�ST�J��y0�o���Ww�c�趥��5�\��m��AC�Y	iHq)  M6�#����7'�"��Q7Zz�3�U,��d7�Qf�N?@�i@���Ƨ�y�g��5�/���,ĺ������σ2|+_�kMU��}��>ܳ�1�^�ᦍ�9���}� �����o��!"�-���76&��(tHc���<o0�y�K�א�S뜾Ƥm<ϩ���:�K2�;��ތ�V�원��2�]ʔ{�=���ks�7Ǥ���Cէ��pO6I_���Q�0B�����?:���"G�΄��&Y�����"��_.cݠ�J�AI��e�3W�+|�Α��~.�h���|�d�G�076՞U���Oy�Gi�F�	�Ҭ�N�"���$<6t��@����8��*�&nm��]���D9�Dv��>�T��e�]^w�
�YT}��,ӊUE�58�/��|��
��#��p��	�ޡQ'Va�;5KF��*�WU�{�Hȧ�1����5�?��^�<��X���3&��Y>;D�ԼF!᯴��i���hT@i�������e�P7�s��[=��g^ ���a-k㷆�LK:�==�4����6�$T����-$�D��f��fށ+.*��@Z�����v�ZR=�|��oc*��r���z��Ƃ��*�t�J�SQ/ã�6�@��ĸ P5��J�}���<)���,[C�I�;�9�����F��iw�wNpu<O��S�T�Oz�U����X,�E��V���I����N���#���Ə����[Ll|�kK�v}X+5(��f1mũ-��v}^!�0��j���(O�o����8��R2㥂�����A��jlb�������ZSvď�'�%��c�o��0T�Q��U;6j{~�������M�����frC���SV�̛��d�)����"8R'1n	�/-@Ub����������@���#��G��' ��)/%rn����?��r,�e�wt��r�8�@V���~*ܚN(���m&�?�87�*	�AVgEM4�ځ���������Z���|2Q����'@6���1�+u A8����3#����2M]���G2� �&d�W}1J�0��#���c�-(�6�����.�H���K������b �m
D����L&���>�`)ҽ=�0QE��� ���:��0T��e�ׁ�[&qބ`F[V�-`��£�"���ߔ�׍�����@�F'���7�4u��Qް`����74&�Z���eJs�N�����D��+�0lc�;w*�)6���	�o�H6[<x�(�7�1�u����Xvs���x�#Q��s�pMU�=��P�;Y����C⧇+�c�i���`�f���A�>6�K=*������������Y�P3sQX�T�w�L�c�i���R���s�u�)�ܚVT�\����M�Eh�iO��k�K��q���h��𜧟d[��L�7{ <�bgV������0���b�[vH��F��&�'��Ͽ�Zv�K�va5܁�:qW��8+��Z��`>a�?z���7���x���qJƖh��&|ǅ�+�i�������3R�Ľ����R�Ҫ�g��;yXT�8�Y�iV0�`�V���{�ʹo#��Zu5��QL^�Pj��o������^F?\�����{X��z�4��*�um��ҋ��哒O�W���Nr,��e�2�wK" �\���v�w����N�[�$մ{�Єi�蔯U3��WXM��j�+D_��i����jJ����>�&¬6 ��Nn�@��<|���=�o�ԇ�[����|sۏ��IxԙEA?R�����8:�nf���ǒw�x�h�G|�N��g0
)r&H�M,doZ�H��nՅ���O����M<^��l��J��3Zr%�����E�o5}T��ݴ�4 YjZ��<��BEr����S1@��{[��?������2��^v��za��>ތ^��1��w��AC5ur�܅n�*c�!�VAHBj#�
x���_�� AK^�w�W�"W���ιc�N\!Q��r�++eF��̇R�<1/<�,LfKR���M\�cF��T��&���TS.�Q5�Au�o�X/1:,�쪣�I�N�e��N^�E�@]U���G�l#�]A"3��Fٙ,h����N�i�?}�Rzh��$i��c����8���'�k��ئ��W��񠌓�K��z^z|���P$(�]�0&�a� �!��hpF|f�͑�X�36�LM�z��I;�9m	���a����H�*c�˘��1� `������%���Y>�fXv����[���l�Z� ����=�"����䑩Q��J��g<�N�'�SI����>w�e���RKnR6Cjz��c3n���ԛ�=tsC^��'~��st�V���Mw���1I�%���sx��~�!ԏ��͋��!��M�=�ِG�.�S��v
+
�����7^�O��}����lt5^D 
�2�hA/i�k�^�4E�&$��u�kl��H�;��S���3eK�-롣i��S�+ޯv���6��9İ�R�ۍT��:�Ev�2�u�c�)�ރ�FW7΃�Y���,�3~�r&G+IQw����JUم5|)��X�
�#�y?���7���S�`��B�2�Ss�ݢlH��	�obb�`�!1G�+�����B�,�)g�c�r��O�V��Y��/�i!=.H�	�������i�6U#�(�R���e��X"�����x�[o%z���.{�r�k��|h�F���=f���W�I���H��i��6_�)�a�a�{�ښɼ���B�ڶ,9���)l筒UuH&齪���	��e�qH~
�a�q̽r�t�)��\P��w��5�` �pJ3�pա������R!J���#��;A}5H.��h5���V�]�i�?O׃�6^ix�Eu ]�(�,/{�l�y����=j�z[��R���at"