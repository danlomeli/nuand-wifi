��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� rā�SZ )����C.��&0C]�-��[�3�-���+��պݣ�k�J�vo`�A�����f����u�X���v�=�а���]Q�Wۿ�߸�=_Q�X����j>��Zw�K��SvX��ƥ.���#�����Z�0���#7{��\S$��@1I�QX~TQ�E��db����۰� ���>0�%�9�j汈��}��1� ��2���h�G��SeY�a���	'<x�p��k�H`�H�j^y�0�s�78+���ֳ�`�R3dW��_��{p[�?$�s0��#�zS�_��bH
�c�p�IL7]� |����Q�� ��Rr���=��E즕2%�����`�^��l�q-�]�p��jf��Ӽ-f%H���ȳ�>��+���M�71��4_�) 3�46h�rb�J�W� k�h~K0�>P$�_n)���5�r�j��W�J&޴o��$>��6��ŀ�;A~<6P��K�~��f��*I
�Z��}`q���ApC��n���g���3��-�іrO�mF���,�$��@�BI�q�}��Ȥ֐����î�䂧��@������U���vU������ �T#K@f�㯁����|95<@���+�-�)�����K���FI�k���*@�m&���
���ma1[�2�u�I�\�U�yu���o�|��2����;�W�W�}P�K>%5�'�8���׫=����k��,�t�M�0�8]q3���Nܺ�^�5Xz��t�l���&��}��ޠ=���< ^�8�$�2���c�=@Y��ɤ�#Z�i���'�*G�����*��2�s�`偞�gM
��㙘&P�<��4���Bj�������8��Q�>�R(g�g&n�80ץ �L��׺��j�i[X���?Hk�K�����	�M�9^�и�D����NWQ�z�^��2qp�KQ%��h,.�Xg}Y���ń�	C�O@#������Q$����[��:9ܺUN��M��pN[�D��G3�G��<U5�d�{��{��3 ��GC��9�w��|]P����t��}p���������ι�!:���~U�'�G���!���=�C����g��Q����wk�aqzɦ����~ޖ�\��2!.��&9-9���{��B���E�*����ƛx)Eg���/��x�H}u�Ws���Y��C��n��~[k��il�L�_�/���7�0ʶ��E�VS �q����G����ws|'HŢ۰������`���(:�˳��EV�X�|�m��o�e�.7Z�\���z,c��y�H����tg���wo��
���,�#W�E�
Jl��!aF%ا����9W��j_%:��[*zO�(�0�����hk��F����ފ)�������~�uws�aY����k7K�a�1������ʸ/g:�3LY�����G(�.�X4�q�	���&״V�uw����|���^�u��wJ4�w�F�YqH�:@��!��K�n�1�K�3����]�8c
N'�I�1�SH��2�)e�1�m'�
�X����z�5W^X><&&X�*��s$�.d�G�/�p� �%��8.��N�t�U�c�ꘪ���M\O�1�"HWF�C�>��$_�u��4�e��6��U}�<F�*G������o#�|9i�S�:mm�y�O�ߜ��zo�fKSy�����gT*���"�5�u�¾%���u�j�����L�r�q���I�k2Pv�Rq�/������
MA��s�mo�ȥLqt�9l �^+M�!�8Ƚ,bF��!����8s��ȡ�QJEy��D�G��d��^�m�݊QJ4��
�v�C�N��ě�n�B
��ے
�5��^ܩ�h�5�p��D�v/y�gc�4`�^�G�|�a$<͚j�v��}�q�(�s^pt~b�s�� F�l�K�xs����[¥����ܣ�C�(�'?b6/��oG�J"�.��I��Η��.��PD������[�� �L�?�$6 ��,d Fd���ZJ�x���D����nw����1�RD#�Uv((5���?��pd/|��1\ڔ�0~.Ei�e?u�i���l)XZK��W��V��g�4�$��=��k�B��9H����XcI����H��Z��0lÜ��Ms��` H���ĵ> <C�-��������¶2n���ѣ�� ��@?�����9�S�ӛs�B����p�N��3��Y��S����$ʗZ�h)�ߌ�����"��1�$����x�/4�{�W���H�6'��&HN/{���4��'gŌd�k���	��g��*�%�PG5��4��|~��ԶC�%XnX���T�~��m�8�\�M57�S7p)�V�{�ut�|1�x��xk�oAeB��x��/��}��fh�^ؾa����8��⮹t/����v�~��\�!���]�a6�uѩ�zp�כ{P�� c+.ԭ�+��W���T�$E�U�IC���8�B�����{EdP���ߧS�{��ȱ�X��'T�e��,tAv{ԝz/YB�HS�](�e����� ���"��=sw�y�%ǽ�#]��q���Vw�'���
e��_�p&�(o�%��HM��X0�~�go����i���ּC.�ڪ� �r 5p�Z�c�J=�T��E���陮WWpE�'�{�!�0ji�	eE9DsꞳ
�	wf���9����u�?JƟ��Z�g�T�hG;��1ꖇC�S��y�˓�W6i��[0���XW`=���QQş���}7n��ę#���d'{�;U �L�n��ԄF�5F�*A�� �F��8�L�	Sx�N[��h(�~r*���YL�aDe���D\=e��&�WP����x+,�	u�B �֝jU���o�� k��i���jAWƛ�t�T�1�����3�%��e�*6�Uv�vڮG����C[@I�[v�l$7��+��\bh�8�}u���*�١�jy���$5�ӛ������5�j�Da�j�jT!��Y�ξ�u(,��B�y�� ��Vڹv�m����38�w7��@�ԣ~Y)�5 D���{��8@=;5fT]�F���%7#��D+�$�C�O���39�akB��~{��%������2�I�ME�M�g]�G��PC�5��I���3)W)s�]��*��"�߅���yx�̿�}4�!��Cf��+:Ў�w�o␣�.fh �{��~O�ݪm�)�Rv����e7�;:��{*����0!��_H���/WE��R&k�	�L��nA�]�Q�W^Ej ��P�oG��ш�*�`��9,Y�����)n�S�]c�� �N!Eg�>��V��u��
|����#r-X�&x��������	�ᖾG�0V���e7^�is'�z�k��[�7�Sci�Eg�1����Q�f�P�'3�����<Oc���l�:�x����'�n"I,0�Z�c��P��*A}��)�2�D�ѧ�߽�Tl8ג�����#�T*2c�
)[��<�������{Wk��<󡬶af͐�Q�N��<�I^4�,�P��b:{!�q���+�M^���S��5��B��b��O�(�a���ƞ�T�B��<�r�ԉ���b��h�W.=��w�5��ڬ�S�L�ƾl(�cu��ؗ�(sLQ3�~�Џ�R�MyQL'�F'�f��n���%�FP�:�qi��R�S�|�ݒ�oa��*�F���׋2Ӄ����ە~@2&�#G���9�R-������Ur�U��Qy �6L��S��!��/�����q,�\|���.�sj У�S�tt�x��b��jHhfj��	n3�?�Ewx���B�3{"N
�m�n ����D�#�Fz7Η��cF���<��ŋ�.�Z��Ҧ{�+p���\���ƽ0و;AYzÿ��ݎH3;jx�ލ�!��E	�KE��I�����i�|1�5��L�ה���D��Gs$���,�)�Jl4�!�	�O|���ekL��H�lw��g$���k�4|�%f0��4����	�9�2D���3�V�f)z�2V��![�CΡx�o�3�kS%�W�W+b�<�?��.F�)C���"���x��''D3A�\���m�3���d��H�Qٔ/��D�I�"����/���3;�T��yro16��~Z��<�{ M`��7!P�vHk��W;x5��tk\�%���>�9O�ء�*8���h��� i���uf��T
���x)�����&3��BY��[]����T�Q3�� ���p�J�<q�`�����?��C�=�JDZ>Y>Y.�m7
,�y�V��ƕʗ:��Fe�������,_�������?��юz^�R!���LA����k��f$r	���ZP�)�#u)j�)����1+Q{�����Y5����TR �K��Rݫ��D�]L�i=�8�B���1�Oa�x�Z�D�X��Y�~+�[B�e��Z/����Lxꚻh ��;V�������X�~
O�������}�@h	M9s�q�m���_��ݶ}��	��d���[T~��+�/��Y�v�%S������%q~ϩ�
����v�H����� *{1�\Ф�D-W`7k��U0�P�~���l ��2�����q�ǒ%����`Ѡ�*�+����5;Zg���ob��{�G����A0۰���Y� �ICu��p�V���lL�PY.AF �'Ʉ���1��@������#D���jɮ�"=== I�Zs^)Ɲ8���w�e��:+gI�M8�!Ul|��/�Ǯ�/8�g6؍�T�������oH\�����G�I�H5��c&^��g��bZ��m'w��=TtP���V��g�A`Ri�L5A�����V�1��*?/�����i����(mM�J�K�0E��7�|��,8�q���D�O�"�)���3\5��An���؉�����p�3|�K$s�S�2��_���m��7z�%6���t�aOQ�t`T2�Ʊ#�[7"���o��(�x�0Wk�2 �<�"@��~*�y���Ma?��bYJ��$�s��=x�����7�<{5��+�E��:@��l��9�D��!�������C�i��|n6d���V<ywۊ:��cG�^7QrOF
I�j��C'I$�k�UV.4(x����0�і�U�A��u|Ą�c,�V@��9�}��սi���w�b}wX��"H?,Z�mV�	/�~. G���%�
Qi2�V_d6Œ�.UE�.���8+�s�5q"Ж�g�{��P<�u������֪��1��W��m���e�')�x�&Q��ӓ!�Xp��܋���9���,5���1kBx�2K�Nm%Pj�� `8:�ė1�or�=<`��AV�T�`������R�@쀘C�p֖�(-��#,��֬��.��.��.z٧� �(e��F?9W :�Ӌ��|��p������|Ȭ��^H����l	��,���7/#�O���変*���)x���i�D��U�P��C5iK�|fiUK���f�Wy�^�5�������F�;�N�rz����	����������s�.�\�\�Fϕ)�L4��Uz���~�dx,9���/.Xb)���_�@X�s9����U�(��ú�숐R�t*|j�	(���lJ'p��v�>4Ұ���,x�0]Wyַ'�	�7�1��hz�Ij���%�k�X�����э��z�U��������^����+~i�����x5��pb���VQ���|��*D`6wI�����E�����>�:Lf/��Eʜ�������Y��+�h�*!�(�+���A���ȹd���� �!�¦)�O���l3{Rpb`[m=��w��1M�1e�QۈQi�i'U���1踤5����:3�k��$�6G
_�N���	z~"�v�������?jė�/"i�{��D�=>V�,�Ĺ�y4`kS"7�G'�ta�(-BJ|� ���^;��l�OǮ�m��#��ސ,j��>�e�`����xt6n;�B�w��An���odc@�N$�����
QJ�A�fDa�~\��RJU����د8+89(��(�C��xZ�����w��w3���^^���
L0�B(ҧD6VZ����"
덕7;�O���띖��NM@���o��e�)ndc�ۓ��)����!��F�\���������Ppc�^�J���?��l����
C�1��[q���T���!�^a���������<P�Җtó�ͽrߵUja��+��?}b��2�I��
/ۭ�#hg����@���C�͛��㤤���$�m������ ��n(6���Y��O���*� `v '�a#�!9]*���D~.�3t�N!���h��%n8'^rR���:P��-�Z�?�D���+��I'<�yjϓ{:�G�_�а���h�*w�#9ŷs���!p��_�A��s�|�W�AG�eI��߳(5o3l�|��'������h��>�k/
��E>{r����Q@=L��Ŕ���ޱ��*g!V�L�Zj6 �����=R�1����3$��[��3w������b�l>d���>N=�"�քE7�r�g���c<Wt��,RGG{�h\�o�x._�4s�I�T�TX�_���
�;�js5�*S��C�͠�6X����<��Et8'^�ڶb֛L��c䧅����#%_U��K������'�7���틵�q<�[�1���B���g�`�N�@P��1T�����t7�g��T�@�c��g�+�5�P�O��̀'�q�'}cg�x(Vʟ��~%�#S}��>����}���dcU���$�H?�V~��J���}C$�o��>�Єk��\�0��R�vvQϥ]�Z�N��Q�^��h���@���{(����M���=\#��r����N�����Ҧ�V��T~�(��obm��/o5�T)�{��[�sV;���(����49��5�X�3g���q���٭��ʺáx��3�n�Q �)F��:��v*hf��<c8!lM�Y��Q�)d�|z-�rZ�r����T]H6�c<M8J�%ѳO
Y�}A�$�}�* �6U�=���Yш�kontΑ����(�dK]N�MU~~�D	��2'C�.���1��.����%��??"$8�	,B��O'��2����Ȇ	��=�0��G�iҘz����j���1(�&��1��U)
^�JSHyAe%Z ��귽�_���C̫�z8�Htz$x+�]���U�E)0A����~W�i�Qv$컵W_�S�/�ɞQFB�Z���Q ���J*�q60�~|z�hW������F����(ћ�JX��3�E1#|�}�E8��_3K �(��:��;+u��������=���P��ud#�.b��]n�7ma�/Q�0��9A=�l�������F��h��%��w�Z����ϵpOl턄r�ߒd�ʧo�����#�vt|n-�9R���W&��C2H�f�����/ڒ�I�@�<���5���|��;yw�4W��j�p�߫�s3��a�Ns߉�