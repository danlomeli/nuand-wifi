��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����xLM�����`,5?p�"���N��}߳�^'��v�Y|'�XR��f����mM�x�p�xV#ڇ��76{��)����L���h�:��+A���9ߨ-� rā�SZ )����C.��&0C]�-��[�3�-���+��պݣ�k�J�vo`�A�����f����u�X���v�=�а���]Q�Wۿ�߸�=_Q�X����j>��Zw�K��SvX��ƥ.���#�����Z�0���#7{��\S$��@1I�QX~TQ�E��db����۰� ���>0�%�9�j汈��}��1� ��2���h�G��SeY�a���	'<x�p��k�H`�H�j^y�0�s�78+���ֳ�`�R3dW��_��{p[�?$�s0��#�zS�_��bH
�c�p�IL7]� |����Q�� ��Rr���=��E즕2%�����`�^��l�q-�]�p��jf��Ӽ-f%H���ȳ�>��+���M�71��4_�) 3�46h�rb�J�W� k�h~K0�>P$�_n)���5�r�j��W�J&޴o��$>��6��ŀ�;A~<6P��K�~��f��*I
�Z��}`q���ApC��n���g���3��-�іrO�mF���,�$��@�BI�q�}��Ȥ֐����î�䂧��@������U���vU������ �T#K@f�㯁����|95<@���+�-�)�����K���FI�k���*@�m&���
���ma1[�2�u�I�\�U�yu���o�|��2����;�W�W�}P�K>%5�'�8���׫=����k��,�t�M�0�8]q3���N���GvZ�i�+ C�e
��Ќ�S�v<%���q��e_��
�k�夞��>ZO7E~��5k�TW Aod��eE���G���ɑ-'���?�G$����ќ����8ɸ+ 5ʗ���l�d��,�J�
�^�3b,�����J����#n�zK����z�&��;|�\�^���'e�W�����">�w*	FO�Δ��v�ƺ����U:��#�����2�U6�vZ�EsYi���h\x�Y��aD��,+d����Z���P��W�L=��a<ѫ�ufK�:��W�2��Z��CX��D�;���x;�H��LJ?�*��	�5�G&�G_�]��d�/����b��kXΤ��+"sY-��ô���!"���EͲI@���c����
�70�`/��O�MWtgǐ��FC���վ컴��J1!���z���j�*5���u�d�zP���4eo6�"�4�ݑgo����l�l��+�}R&�z^���R�"X�����@>�O����V���~��>��2���|�2�Ѣtn%���s�c�1K����z�$�slëL��^>�ˀs2%�x�]����J�b6a�C��Ìg��'��l.�@	Է��p�c0��Du�4"���vx�������Yܤot�I32ĵ*�*�O���8��ګߏ�~���&�Px^�8�UM����lp�Ы"0]H��8�6g�ݽ��Q8y;�Er)1X�Mc.�]e��2~TlZ/�[��o�ohH�e�B���j����0xB���5.��3A��ԍ;Rq�W!�ω�-�X'�]k�irHN3������j���ė�����\,��RP/FW�+u�Ύ���
�� ��1nW ��V�:~��d�;{Y�v uH�8%BT;���N%(֍3��W_Z�<|�0�7!W|�-8~V�b��@��W�: ����0��W�y4���V�����KĶr�N\
�e;âĩx hFҗ���Dѱ>b��pf��.-��V���,\�� >6_��M�.Ҳ&�~�H���I�k�Ġ$�"������[w��!���UD��ZEү)���<x���C���?]z�}�.���N��)�|&I�{v�D�n&��������68OBEQ�Q��7�Ax��'a��uϬ��L�i��BB�)���.���?Fg|�^S/�\R��[V�W2�pA',�ഘŲ����b`KA��b����靹���f�q��)抳�Z��L����cv��^��Ԩ|�g��U��>4N��� ���k��T�<�Vh��	M,}8 "X�FҌ�[�^�A�)aB�� �	��r�}y!�ɏ4?!��exa���zo�"	UUM��,��=��?��m
��}�k����a,��xV��p���+�(�J�ػ����T�/��l�N(�Ps�
�	����CQ�8o��FX�Z�P	=�R_�6�n T�FT�62�i��ӹ�t��ޞ��i��
�N�@�֍�}\�n鼺]~����el�;�c+X�	`n٬�p/.L��:l��$)�,�^��H 9�D�K`d{�S��������}�]��������׾f�30e��(�r]���qtб-���e������Y�w���᪠���#�~w;��r�,|χاP2���*]�jn��3I�(O��{�9Y5��c��7����
�Vc�[e��?b�2��L���ׂ�B�BM��_�=Q[(M84H2f����W�C_�HP޶dHM�2@-@�K� h��,͊h�0@ɾxi�S�"Ր$����	�F��3�%�Tp)�R��v��5"iM��;�9��+n��z|_�d!��ܫK��L�)����/�hH�
�Q;AX����v��Oe�n�x.y`�[�tbژ5Bc��E��0֮a��?p��26�gj<I��nU�7/߲�J@����9:̭�.B3��
g[t�;s��:&����O)�[C[�l)v�����e1���d���&s�"1��b�Z��pz� �ǀ&2"���YE1�@t=�g��˵`v�B�|9�.V�U�9�Ń�tYg1OP��0��87�@�$�&�*����g�}�>�N8ԟ2�ݚ�sPL�6)�� D|���'�|�u�j��u�iv�JuZI�4��N�Z����EU��Cd���e���ɇ�Z�aL;�N2�b?9��T�L�S�Y��MIo�`9m�6Yx<��9�)zE�E���Y��hV��](7�%�����M�~*�O�D�NqP�<����~n�ύ�c�e�Y��gǱ	���K��J���n�n����t����(�p�π�E�݈e�7��.���)5tz괕Bh�lQ���[���I��J�@m�B����t�S��k<���=�]����J�p�­q�T&�M<��0��s��?��ۉ/���{<ɋ���Ӝ�t�V\JbA��B~p)O~����c�?�Ӻa�>b�R}*�D�_��9+����ai�fH����� �v�y��f��.g<)O�4]��2�H�;����=�����3k���u�*����b�خ�j|)�`qg��0_���Q�u��:'�<Dz�T�+Uq���#�L�.�vN��ErA� @����e[p�^�$:`N�r�����m� �x:��f���r��X�ƿb�@-]��U���Q�%��ĦSn���:h���e֦_��Θ�y�J�4�fX�4�\-E�nRwхUwTOPLp+�	We�4�w�0�2S�w��^r�K�?�_]��3۔;�Dt��^ʄ)�*_�n����=�Z�8$�#���<�����OA=+pE�j��X��lT`����,av��B�R�mH�
x�;\���()����q��u����G�<�/`�`��ط�z�t�"�����Z����xv��^*k�Wt���!�.��fxg�e��~�qiQ]���#�,��ώ	5m�^or���"���&��:}Z�� �3vh)�:���X�M��y�P�l;�Q���g^*�.���Zr�]�o~g`(|e1.����p��ZB׶��B\����}j�#L��T3����;��u�+�O�)ܐ���|���$>P�W�K$v11���1Gŷ�aU�c۱���Z���C� �ɬ�t�+�:6��� ��Ӡӛ��e&�܅ftۮ�U���xV����O�>���y<��A��SOL�0o�̹�Q���"�d��+llr�c�8~��*ˣn򚙘i7O	h-=�0�v���q$φ=ňB�HW:���-�z���[�(�t	��#1��ZC_���0@1���V�s뱬CNx�k>6�����3�0�?��8���k^z�g(M	p�PJ�U%�m��O�֭Z�Q��(E]5�	 \sX2����6�p>	qF���Y˭n�Zq���E4ה�t��`j�N�]A�!�!�ԦϨ���5�Ps^�7Iȧе�����=�r
���V��N`+iG��{�� \�un�v��{h�Z�EO�������Ä�l�|��E���<.��?�{���m��N� D>a;����� �8��<_w��qBK0�L�u��N��1��Y�)K3	�%�n�5xi� �� �
�OP
����ܞe;A[��_�=�7���������6yi.�92�*�nO��/�ݑ_5 �1�k�I2��&���������ĕ���3.�h]��i����;��r�����'�]hK_I���{�(��dY�����E2���7��+#����jpo�"IpxN��J�F�}�g�#ޞYÕ������
���٤�4�1`��#�a͘�|�i�����f����tmDY!bba�lĘ��/^&�@���Ip*����V	rk!g���-��5�#(_�8��v��w��7Zg� ������;ڱ�Q�9�;�ÜP�c��Xs�Z��d��#a�_����Ǚ�����k������e��Y����nE��#�F�d ��}w}������h�ޝ]%=�sDhŘW
���ª�_�A#��r�>���7i�1�c?$Ίvx^��v³�;w��u���ql i��xW�K��u��T��B���r��Nc�~�޷��֝T,n{�6k�9���#�� ��L���Sp�`�c��Ki{s�!�aE��k��<Kw��y��$ʹvu����]�0�[�N��������F4��6ɯW�F����ƾ仢 S�ڎ(���H���"��R`�p`-LWո��1|%h\+�t����Ux�VC�4�;�a�w�'-�Q�(A��[ٜ�����J�w�^uխ]�q�K0�����B��^��"z�T��!���T-]�J�Ȯ�X!�5�xT�
��-px��5�G�k���lr�U�Y}�Y��Jio��ˊ$��=�2h��n�FL'�oM^:ºB���a�f刺�gb���V�?O�����d ��AW��bS����<o����Rx�:�>��"��s�4���>}�R8���&����LW$�x��3�K3�}��Bi�����0�|��*�Ѓ�38�x�:�$����Ӯ�vэ>�L���D5���K�Z�E��^�9`Ʊ)�H-m~~EF�7�-�hd!�bBH��ɾ 0��`C�.D��G���$OX"U�N����ğ��X�z��8�$壜 �Ơ/�r��>�"]b�"�a�Ch��d�n�5�C����.��Y�2��وd��S�ZT�������A-}�%r?:^�ע�Z�$�x-i�aP��t��M�F+����&���c�sD���[`��P����Y�����J9E`�FFp��p� `݉��C�`��%��"/@w�d�+��d����^�W�6�_��r�Kԇ�ٔ�y2�	��JE��}@B��� ������_d&��m�� isǥS��c^e)���S]'|y�f��Q�tn�B0��D�͓�k�4�uÜ��wu����lxU�դv�3�}�����s�P�
=��-H��G���}�C�O�%�{lz�hI>{p�g��mCX���' ��\|r�ܠI|��xB�(G�hY{L��=S�����br��k�ՠc([w)��ԨC0q��Ģ�3�=B0K��o%���M\�:�|����LP��{R��}W����(�G�ٽ���)�{�p�M����D���őݧ��wunt�LD4 U�p<���
IfB-�/�z�y��}�4Pw����8V�%�_��:`TIS9�'F��r#�y�Վ��x�H���B���i
��iw�H���1��<�mޠ�ǛЊ��o-cR9�h]���W�[����Mi
� ����wb���+�oA��Dru�b�9W�{K��<t���B�HqT�:=#+ �I}���9W���Y��� ���ɝŜ}�(�@��`t�O����������(}+"a�UI��a7/7�@&=O=Ѭ��\��x9-O�u��%Q;Y��>���7b��G~�-���'� �jO+���+X����6l�3l��b��+@�7�3vs��r�3���	�hm���#%]�lnT<�1�:�w��Q���o4і+Oj�N0�q|�m��8>�/�ƁB�}Z���^�:`?�!e�g��m	��d�E��#�
]P��RC����W�e��p��s�����/G��Jx�ް����u�]����:�$�����5�$���힭��9����i^mm��m��܁��^Ul��2���x47`���ݹi>�!���8z�w8@����0�!�w�0�}YU�$�H3�i��}�a�!%��	�4p�Xn(5<r��//�-���ޮ N+���4��G�5�0��"�l*�C�a~���;.J��<�+a���H��[h���#�Ƀ���.�eJ�#�|e1CB�݋uy�[<g����_�w�"{hطM�
B/`Hr �S+�_w�"R�Z7�9��a��
w���:G�-�������T�+�Hs��e�{����u��@D��Dq�e'�f7%���ߕ舲3����ȹa���X�������S֏���z�}��3n��7���YZ������)�������j�$[�	�؊�A����O@��QJc�$��}+�:;��]�I/�HS��c�􍬩A�^\$
P��.�Ѽ���:��χ�ۂ鼎�s��CU���������j�&���TBp�*�>S�T�$`��y�P���5��YqS�br��/d����m�Jv��o�;���Z��c�w�%�����mJ3�>�iX���O��g�u�f�m|���#ҡ�;Q\(�pI�'$ƹOX	��W�? ���V�����q[b|�<���Z�q�mM��P�Q/#v{����=�/85��F�b2�V���,�Z��CSyJͶiJ]�@����#�On���1����ܛ	;#�$����Й5�+qQÜ�2h��^����Y;̓�:߆�A���b:��,��Yo���}R�	�c�+\��Z�z��1$��O�P��$Vk��RDM��>A��X������ص�������g	�l���qTү�>�u��UQB�uML�V �������R���0&����e���IqwԳH��E9y��Imw����E����yB	%����s�$PV��6V�Lk���V$�����H>�٩�َ��V4V�8w�ϻP�y}�)'"��W��!O:Eɕ� �V�f��d
���:D��t� �����	��%;�ՈU^��3�Yz-�����}���(]��3V7��cf�y�����עx���9Z+a�`D��;�I�F� �i���;�7�;7K���3��w�}9w�UY�v�v@p�$!��z^g���
����Q�:�*�����?���j�&�����k,	�l��oE��1p�{Fxz�`�?	T�"z�g7�q�^��ϗPa�Y���0˸%o^�(��[%fs��Nnj�֪HZ([���2��<������)[�{�W9�w����ɻ�J��2D���ʎ�D�;�̷b���Oyh�֖w�@��w�C�7=x�F7�+k��3C��%��cFm�OD���R|4�B1ῆ��5� ݄����ܖ^��OR��lB]`�S[� f�d�mGPS
\p&���}��ԩʳ\# an~�{}�����R�~���"����ut'k$x�U�q�
V=��ޕ���KMF�L����T��'�[�m&D.Pc�V��=:Ӱ�l��@��O�%���t�A �s��m�8x��d9O!��x H��z�FY��`ˌ�/��wn��č��Y�e���/m�[�����*����ݷ쯞��M�|���^�a&RG���7%�h(3�<	�S�c�ӌ8v��y��@��W��*x䪈ΎtN��JpY�o����l�@@NpzT\�=ޢ_qՆ��k�?P\�Zj�ӳ��`V�����G�ً������
M���Qod��!�l�=��h�W�{_������5\+^q�Bq�]|����`"h�%��f���*%�/;s��u�"t���$r�?G!é lݭ��y;�ȢQ�@�{+gh��ouB����I?o����K�S@v},�]7�a�������HQw���s�e!����h�w����`H���%+Ӳ+��t�r�)X�W��Q��΅N���b6�L�P��G[���#�'�,��s�$>3��EV$�|�,;1'���ϙ+^�&p\�=�� �3A�9�kt�A{Ihe6%��C���&;T�淡Bj����&��:��P�`��J�ö����ZRϝ�(�g]U�h��dp�q�[9���,h86�Y�e�\���}'�%��(��35�cYP8���W�tu�I��Yֶ�P���t�l�s�A�B�|�OD��Ѵ��11�����♄�g��`�@];�h��"ß��{-V�S�8�ȹZ�!נp�������(���>j��/1�������y�׫I��C�=�.2ɲ�+8�k.���/�iwu�*��%�=���_��k�����0P"��ǬNcib&�����~e`|^�LM�7
^�k|؈���jAQϑ�f�4�#ߟ�<�!�t��j�|O��];�Uh��v��Q
vi��x�{�6t�q�Y6"q]#�_g��lKm���I{Fв����H�D�DT�i��3�+�^|\S��-�A.`9��y���|�W�O!�l�����;�g����^5l�0xy�Z]VWŜb�ĺe~�����Ǿ� ر��z.	�76*F���ɷE���ALN����a��L?W�u�����h�:z֮0��B���*��?�ш"A�Xw�G�?\H�H?�T�ٻqb�x"�$q�J��:{q&�W�ʟk�u���9�~��^T��}ʝ�^ �@d��HveC	�[�6��[���K���q�Rb6D���'��ǚ[��?���� ٵ��P���Aڸ+oAj�WR$��@�7�Ќ����i&F�Q\Z?/v���W�1<�e����t�01����23
E�Q{��	6��h�n�'�`�����^���&wuL���\���֐	�=覯x�[�'��c��9�R)Gm����]9t㣋��g�t���˩s�
�rߎ������:��^�Z0P%����ߢ�����I�+�M��h��&�h��T����������"�qp��R�.���w/R�@����/�edW��|f�g7�&��&aÃ��&���+�-�Pf�zq���t����V�~d��4�!B:�uM��| ]e���ԛ��|z1#�^��_�>v���"���	Do;��;7�m��� -�P�]|�GU}�oq ~^�U�Q��#W�I<�ۍ0ō��������f�Q���v���V���(���8輋H	P�z�u�uR��A����{�P}��b�-8�&`搼:^m�H���/c��������Z�WA�Q �ܵ4^�!��"�`O��w�e����(ILcE�K�N�
 �(<��I�"n@
�!�[��{.0x+�&3\���@���HF�����8c���o�:c\�>mT�j��1���-�pN�Ԕ�I����Zw:"5��Xrzٜ�4:�˨�f�bvhݟ���A�אcJ��|"NH��SQ��9k0��E�U�0�)54*�h�i0�vjP¯�Y�Y8=�e���?���y�T��6	�ޫ͂�b���k��m�w����j��,\5!��v�9�y��p�wX)�UP{�5��܌�Z��T?	W.$�@d(սv�ʑvv:�ǀ�&�.��8\��Ko]�n�C�����~�y4���g��"����3��'?.�R�V��t
Xv�f�+�����z�B��a�0���2���//~en=���{��(���mǘ#�����H�dD/и!K?ğWM�L��)&:�׍X��EQ�Zd1��O�� �ߝ���!��A�tܟ,�@�-���9V�.�i�9?�C�N>�UbH}*��8,��ף�z#�����Msz�
�9�^8]��Ղe�f��JVOr�7g��h�o�n�@�5s����'f�xW!�،'g�V�q>mQ�(h_@����pK���橔��Uh�����!;�5m�f�����k��~B�@���.�URp�>���b�6�Jj��.� |Me�C��W��!85�4�z��_��6k���H��]�Ī��.�����>Q�O�����.������9)q�+���|m�.�I�O�*�m�&ב��Ѵ<��[g�e���ˬo��2�׎u�y���Rtg�|��!��	�z��IO{�h<v�#l�����,X�:�X嬖�yxB�M埂:�-iӿ^?=(S	c���S/�T���0im���TB�ŵ��Y�M��t*�PW�|W�I5Q%64��JW��N��k�\�4��|Y�j̯]eLE�zE�Uzl�s���CEh;�*0rl���a��%(��ȁKWs��Y#����|��cg�d;�O�$����GG�L��y.{E�qG���
�q*cJ]�1�OK7�R��p����ƁMw�*��H6C�9�%�#e�;I��I#�u��2��Q$_Yt��ʸ���իV[�@������ EH�|v�����e���Q՘�����uh�����f�zD(�ח�	A_p-�T��"L_]"�&3c�pay����o�����Ķ��r��@���bPuC���]ʾ��;l�g �A��n4
�}ߤ�����K���U�sܱK�o�:V0��gh��rf�u�����f!�Q���%�{x~��{Cu�������4ęB'�U����BZ
�����Ou�7MX��d�t�h�G���+G:�(vYS�cE�Qf���J������c7�^�b���wP�g�'���k��L<~��@�O�i\ ��U_�m���/*��,ۼ	�0��pD"��Ӈ�9
g��О����J~��v��ܾ�:�(����] q�V�!�!@^Y���J�ok��Z �p�a�0C0%H��}�����g�$�۞t%Ց�j�N��}�Yk���}M܋k���qcf��x���Vy�����\R��Oj�6�_։4)n�޹�?�����6�i^᫛t��I��TpPRP�I��%�&�q�p���g�&7ɜ�5�Yb��	�ߋm�����nE�GX"��bVp7_qUCb�4O�(H��8�q8�z�jP��	�3�g���c��7���=u�U�ZH��!V����R�%�ԗث�F�/'Q��hNF����M�n�����w-�%Wid
	�[�Z��r���yh~�B����m�E7}�7x���j{-�MOL3��(s=�a'9:f=_�Йף_)"����֨��E��oi��ƌ�M�%�^������*�Qۂ�[ ��O&}S��L���&:y|2��}�J)�7Q�8���]��E �,���⼐��tX��t�n���ì5 s0��>u}(�W���uL����4�ݾ����蘝��L�K�pr֞@����)�n�"���	�O�7{V�c`O�n�v�]zv��g�5�5N������
7ן �c�Q��E���g�~?AE��-��[I�E��u�	���z���a�{6B�ߥ4���>9�.A����?th�t�>���G�ּ����iR��ǉm^0F��i%�
��tn�f�#����XˇW��ɇ�?E}�-��ƫ-]��n�� .%�s�K����7x�'suj^>���$����X�R;��82�� �C��#��m;����H\���*^��33�Jqo����	s�r߾�*����'i�u�h`î�%O0h˅�Wc�N�ФLi�,N��sȻ�5�>���ujO��ӊn���,�<b9�k��x���=X�pje����rSf�H��D��UNE(������t��$����g��]�<6����WoC�[#v�)E�cUC�jɌ_a׹S�D�eH�^9�P���iu�����w�v68��37b� ����?n��|��"p]
��T��|o�jTo5��� P�殺�iMj��=�e@^�2�\�������I˹i�������j���p�L_��3m-���}�j��T�	4��KFl���nSV�DUV�-v+ �e^�bH�>��^���ǚ3��s)��_>�'M7\p@��K4b�E�PR���j$~>���FF@P�}-b��p4k���߱��GG�
��W�1,oCO�zf`���6����!�p�nWcA�����B���ĩ>8��>����؎�(�_6�Q\�KR������wzAS3�/U.!��i&��U��&ddA4�WK��Ƥ��Rl@�jJ��n
>��]�[a��H� Z���e�H������m���-���G�V7`a0�����l���r*<!.�� )���yF���8��9ٵ�9e������0��>���W��]"a����V��?8Q�^��$]�Yd��^� �]�WUs	��#�8�����_��B���V��Hw�>���k>G��Kx)���^�~��LQp(�<��X��ĊlNR�0H�#�q���B����m�=x!��;lŝͽӱ�9d���m	1SJ"(�?�2$Ť	O`����0���4��Ot�
 �&Aoi�]���,T�����(QYa��b�/�t�z�4G���馡Xw�q�Eo���<��%鞸s��Y[��_�|���.�IT��p��ag��L2�\9S��m���%g\p�pVT4���4�<�qg�e�)�b�I8��n���m���wq!��3��М @� �j�[>�f���7���Fb^����V>IJ�{$�xV���~���Q���}�ص�F���$����l7-&�G�+���xX��Q�G4wvk��mi�?�Z�!Rh����O��	L��.O�U]�i��J� ��/w���j���G����-�l�3b��4a��＆���B��B�`T�W\�wmt)� ��8�AY�8���#��^y�̣���&O&�ᑶHv	\JIj�wҡY=��PZ�:��ڱ��L�V�$u�w�X0ۥ�(�o7�c2���h5�*la8����ZA�-�O��Ƭ��@��g��=|���
�T�n]0��Rqw��=F�=u�x��+����Z��$���9CD��� ��f;;9�����2�P�}E� �9��1w"�=�Ɖ��TO���=7�H��k�r��w|�J#P����֮�j���+C�V�"e}k6>�y�ί1xYʑu=�v	#e��901��i��C�5���\�2�+5�ix�1��%Y��EV��K�"��D	�~e���J�нÞl+�ho�Z����Fl�6Dr���QZ��0�Ṗ�^�#�0�b^N���%u����TU�A��$�a"U�V�H�q���t�W���em��$�y ��Zin�eF����H��<l@Q��,����<�l��0P��+�#��˓X0eT�j���)�.�|��ى�,��.�Y�����0�?.�Wr�N�r����4Q�N�Hu���U/�,�3;�z{J�MN1Y��-\�w-IKӁ���?���?�튊���t)�e*�8S���*g�0l�cLV�a!���/�y��Pq-����˷JBq�	�)I������j4b:2�F�5�Y�A��?�A�:��a�G;�1��L#HD#����:"0 ��$�@��2�n��"��+�G۽��d��N��g@�P���.j���lηHD�WO�c��ŋ�=���셮L�7�k�"8j��Q/e;����z����z4���׫������:�}���{o�`5�|��D��'!���+cqL�KV{5�<�U�ݪ�����P�>ܦܤ#K�R �ș������(�E��Z3�_(h�#���6�L�����z��db���+<�՘¡�2-2~�iY���9��zTK��Y�6y�!�^����M�龍F��5�מ������Љ�\&���ܮ��%�ɇ��W�/�f�V��
�~*�R&V����S_w��f�$���\�$��a�4D���ɡ���f�	X�jPc�X[7'��7�I�������jzT��Ư˞��@��)5C�,&���=q"�J@�Xf�U��ڀQ4o��3Kϱ:rA! �r���'�`�|xSڐca9�Vt�"�*�����D����
�bC��y�O��p�����X]���}����v���E8���*�\;�)�5��3���M ��|���?`)��W�����c�r��Icb�q~}� ���F�'���5	sP_� �l�-w$��o���8(2��j���Sz>X�:�k2��*y�Q�(� ��ϼi/��9W��6�wܸb� x�ަqɧ���A޷�Iaw�^<P�ޕMJ�.5�N Y�2��m@k!(�_pW�������
�;���A ����1�X�
�~�4!oN��q$�����7�4��xeY*:�����:�y�RB��cñ}{ɑ�Q �yo�bo(q�x�4�K��ђ��,ˈE�}�1d����a����� :c/�mE�l���	#�[�����7���T��+�6E"@w]���K�����.E_���8�fH�u�Y�����s�Jv���9�`�y�*aa(5��veOZ�7�����ó�>s�C���ǉ.ܝ��ْ��)�/���ӯ����W�����p�C�#z>t�����	�o����w&�4RAv/�s?h��(j]����:�,�n�d�7��դ�e��p|��$��N�?�;�{�j��s����(n$<�����	�e��^���]�s���W�7���Vp�g魑Z4�����dw���Ң:K�qs���j%�[���|��"����K��}�� >O�$���M�c�>b�ӽ�/�JDc�*�U�T������1�iw��p��ҘK3�f�f嘊�Gx_�n��oxRD�O|oęD�Yk��	��/ ٷ�WO�	j���S��	�w$r[�So�^(�x�,똹K�����pJ�N:Ѭy���k��uF.hL$~��ek�4z�٧�V�I��P(�-|isK�e͵��W�Zv�������/W,�@�Br\Z��ny�,W� �ɀ�!A)6*�p���O_�mTz_/V�/aѸr¶�X�U_��H�l��,�NQ@����3J��,��� �~iT~�wj#�L��v=��=?t�a�I���}HB�B�����������G8�)��� 
��&�pV|��g���p���Fm���z��춒�=S�� =�;MZ��j�D���� <ɬ������7�b.���,���O�Bc�ՅKU:|�r��Gͷ��R;�5�ʠV�埌���Brd�<itahJ��.*�t��#�������YJ^$��"�v���Tf�����#�T�gB���n8	�Ȑ&@D��68e9z_ S�u�ח�+	j���-@������K�|mR@v�0WC���Ȟ�'�9��蹬ע٤c���Da�`>틸@B�n�-�)g��S��';��֚֯�����j�R�����ː�W3�Fn�^����K��;� E�7\U�yU���"̀���rw3��-��ۥ�/6�_u:Q�k4�g�(������_���Y��p=�4��1T6�ʏ��A����E�ף��ݝ�D�J�^U����'r���H�3��vk--����3�x���S� Un8y��ͤ��b�+��S���D�u���^�/S����)i�^��)m�~R�ʯ34�X]�&�5z�HX ݌�l�f�(�U<s�5�rX�|-`L�������pM�]{��K��Vo�ʩ�@K��^�J�?��δp���>؏OE�0�KޯdH�r_ˮf+�A� �Q��Q ErR;����V��܇GS����p�87Q���*^%�<�Ѣ�,��pJ�$�]����ίj�4h�N��̭5�`�P�E�w�V}_hI�\���G���a�]�<G-����S��r��,��D����Q���'�{��b'����0�s�9�f U���.�5�b$��"����e ����"����nf;����<�<���)�؈�aR��P��^d8!�P��b�
xNj�~J7@xW@\=M�J��e��=������J¸f�A#�tJ f�h.�cnlw�C�x�l�Ƣ[?IuDycb�?�� �N���a��>�xjx�@�Ǘ.p�	Qi���0��������vb��V,���ћ5w��r�u�O� I)cq���}�}��]�*��#������e!v�ľ/�b �Qz	�F���8�{V��8��:b��������0D��b��-|b������ٹ:��[�H&�9��3���;�������Ӿm� �de�!�Q��%��t��˼�q�j�.����.sjv%�]�隐�
��n��J)4�V��P��'HQ3��n(@ҧ�Y6���ڇ@�_�)p
�=�Y��Qٴ�/��+�i�^OdR?kG鹣h��.�����ӭ���$!X;2�J�]�;7�S�^ܳ�J�j0�:��h�fծ#�ʴa2:������֑N�`QR۩I��kxq�w�+`?Y�-25F��gBp����e��"&��3p ���a���c�^��9�Fcl>éxe�+�Ұ]�P�6�Q�������Pze�Oe��s�D5F�z��V�߸O̀�[*x�A�Γ|��X�c9�B�hF���Q�0��5�˕�13�J֚��X�j�{xp�pHA{~���!��
����f�u��T�ZfK@Ĳ�g
�1Ò�S"�'�K5�$x"��������D�*�}g�a.���8Q�΄�$o\G�Z�?Rq���ƫ��p��ZVU�%�?�p.�<5}���=3��F��>�..z�3Eи�[��.SVh|���B��Rm6�_Bf�P��d2�Mt��sĩF2�=�V�,��X��YmQ3�-g_{��;��OgGW��|�-��|��s��*?�;�kl��-S�}�w2G�f[���4N�t��*�߇��D`!��r�ݧ�i��Q�����/h���ҷ?SdK����2SA�`��Hz��[�{��x4�<G8)^��_�a~���l}��D��iɷR��Ɖ�;X(:��ߏGg�'1�?�(�T�y��l���f�}�Yf���0k)�|�R#�~[%=��?ֲYU%�ZG�^�	���VqV�fxST�~0���V���E6�ۡ$Fi�υ�P�"FC3h|q��Y�M��4}�`1(��f�e�k(%d���<�кTi��&��t���P��4�[ӯuB�h#� ��g^�G;�~x�{K��ܢ_4�'�崊D1��0a��xa"4h�o*�jn ���yRsxB~Ҡ�|�h�g7`���إ���l������뱂��ƞ;>���Z�����X�b����A+P�0�S��T��(n�7�Q^_��Oj��ak�cZ�8&`�S#�5��l7hQE�;���K�q��?R�O�(h�=�I������d�	=[T�F���=��d*���M�4^Oj��I=nXc�/<�u6�N���F��S�:U0<M��ׂI����\�G��.�����^_/ PG1q�7��?�*����W%��|+��xyWKt���_N�# ZJ�G��<Y�(���3��!���-�b����%L��:�k�~�e�\�4e��pC1��8�1��3L����)�߸��?e���q�|��Я�pG��Zd�<y��q'��L��[*�6���'�ʩ}���u���=}v����d����� ����l��nbF��^��G����o��"bُ����zQvY� 
�=?~���xLS�I�i�9��[��CzϴB�OzP�I�i��Q攚PCrg�L.:��<��"vӭ�%탶�jVD��}dBז��4%}bF�1�����}=N:�z#l�垦��؅?)DӰ�{��+�=Q��1oI8��4��:�g�x�];qe-����y�ӷ�M)���~hd*���JWf����Np#�N}!�(�(>�TUAm��_�V8y�@���C�l̠Ŏ��Gj\�����e�q�ej�i�0�S9��M��Sj��cYs�F|�����s
���ˇ�XcPϠ��O�;������k�c���ܒŊf���o�7'�'	s6��+�߃K+����gr������ ��3 	��kS�r^3'�󻴻��M�Qˎ1p�S:�q�1h�̀}��}'��iT�#���Lܢ�I���ͽu5)���`���5��4r5Ӓ<_�̧��Q��gL�q���d1��.}���ک.�̞���ϔӪ�ʡ�ݽ8V�TP
��0���Î��������U�ZqN۷0�����i��ۘg9Jƹ`(Ayޕ֗7!��_�+��'�m�7���L_f����˼~,{G|�}>�3�6�<���W�U\0�g�t-EA��5��
��h�ͻ�ͅ���fM�A��!�����L󘩛}Q>��-��=B��.��֎��o]F<s,ڝ�.brv��Eu ����^�X��k��MZ	NX�Ƹc��xY$�L��/� >�H���)װ�4N�ȸTr��i:7�/��'�c��۵>��y�z�#�%�6�vM�k3�Q���8�>N ��`zy�5��?ʫ|�p�lX~�ӟ�Μ��Źʵ�-���Ӫ��R&���?9��9�)A=��������z�zV��;�|撜�H�u�L�u�g���-��s=]��"��g����(�U	�ܖ\�.6i²�<�й��\:nb��*z�@�u�����GTF�|4�j"�dOd�L[��9����u����R�X�Z���$��aoɬ2��\��a���� n>����^�^^���@�Qa2�(����踞�־	(ۀc1V.+�I�y>NzI�-ި
�f�'%}�����҆�Rb^�D!>���u�!�(�okV��u����Z�?gQF�ccv6;᧟ѥ� `I��Z-���F��!ۿ���Iqz�N#�9��5�;,k.>�~�~��O�.�.��˜��[zTU��_�pƟ�B�N���ß'�J��쭳�_����`k�f�����!�0��O)��{4�Kd9�����]L�M�=Fͥ�������-H����?�6�BE���ܵ��R����¸�?�g��en�ɀ^霄4��!�gԲ�*<@������7��%h^;s�H'*�Z3�v�,���\�QE���gu�`�rz�8��#�j�*�#�)aV��p�8�f��j�h43E�Pbm0��p��4� �%.��3w�_*��Sm[28(��g�����&�[�B�i���lȊ��I����_j������2�4���0W�����J���]�������
i*��������xT��S�v�F�c"sѶ"�=�#6�a3SbM�H��u(���q�9�e2�9���m�M��5�Ez����S�G)���wRWڣ��9�&�Q���:�rA�$Z���N���"�
W�QWu~�$�O+ST4�_[��;�B;����o�j5/x��
D���Cc���4i:�� 3�uQ�:���٩�H}IumT��O�>�����!��@�ڎJ������$M���A�0qd	�\*f��]ouϷQo��G��iԻ�.��'�Yޭ� 2��Mń�ې�׿?�J��|s_���J�mJ�NY&��uo%��K-�Vәh}����>c�aTtv����NH��h=�
�68bH�v����Q����[������ܭ[Y�S�f�7��ߡ�����f@Sp���D(��t�E�z|��:MW��`�angSBpy��N~����z�{�*'R�9^�B��&�m�j�=�,<*��� � �mn{���U�KO�+� ���-�� A�Jea$�t��CՓ�ǁ��ʌk��J˾v,&-�Ck�zǺ]FK��9q]u��%AK���Z�gA=����Đ �Js0��y�Fm��>g��������إ��%/��t+̦r��*a�|�A0a�_��d�d咭�v���Z�䬼ĊU�%� [9p\�}�?O�e��$-��1�I��,N&şϖ#,|���K��?sc&k���Vk����B1�D*u#9�MD�LW+��8�x0��P����$�zw<o�L\&GD�v�m�h쳼b'�#72�4����!RS~62���V���['��Ui�}G�(: �s6)�U`�mI�cQv��M���V~�W�Yy'��AOm�ʽ)�����Pk�j@iZP���CA5���1��}���FYUj���@`���^۲g�����w$�K�@ծ#��	&X36�f����]nU#/Vm����̭���@i�&17v��W���A4vbD*��'����T�O�"�i�YH��ѿ��(��w�
��r���Y�=��y��x�>��u6l���sg�*������{��v_�z/�+(���k?��?��4��b��0t��f���y =�"	T|�-e y9�6TП��V<~hQ���*�Em���bȺ��Ժ!��j�R��r2sO���,&#v
XM�0w���p-�Ñ��M�BP�8��~@��w#ׂ+V�ߟeR���@C��x��b���M^�Z\3�8��#]���U�^Tę�⢽*^V'�"�g}F��b�nH�u���W)�-�!�P	�V=hfwg�t��o�d��K�)ٞ{N�ǰ�ܴ���̆V��ƛZ)��اC�GCA��aH|uRU��b�OC\����Ĵ�g�G�Q2;'���y}(()�x���1>�H��4�YЅ���K�<�J�:�ޞ	��7NH���e������"^�@f¶��z�~*���\��*M��ڗ�m��<���Nt�2���9O�S)�<��$�����F}S�����Ett;���E�*��1�)�&�=�'�0�������������!hA{퍬Q�ݷ����(ZV(@1�d?���f��mZ��Mߧl�z�d���;<�e~9f�A|~�o��l ��)�w^�
up |w�M��7~�>b,���T3���~�=�J��䫇�"�k)�
�	Q��;��<b04��pSo
 Λ�55�Q���Me�W�i2�A�|z�9��c;Nق.	v��66���%��=�HzL��=6���;`����C�c!�8�ikes���"$�@� ���r'mݖB1�/\̚���@�0��a8�j���#l�O���"A`�G��7�wM��Xt!�|OY8.�^ɂ{C��.?�~q{��:�X�}��P�)&��)�EϞ[4�R��&� .2(�=
T�����7G���ˡe6�Q	)B��p�y���5g�3�Ĕ����?A��\5<ޘŘ�V���!?���� ?'2MU��153�r��2�|��jO��ݵ7>j�bj-c�5�3��&���rB�#�'EXD�������<�w�9�8Cp|��+�͉� ���q���C����[k(97��
{�5M{��[3��7�Bݪ��lp��*/�M[ٽƗ[X��k��	xLj�rk��nQ���1�oy�!���i�p�.Z���*|�4i�Tz]��Ⱥ3g��=��x+� ��<Q�!���L���5��P\IV��W[|�?t��g��usB�lCv��Y$�ƃ4��Z�Lc��������\��F���|':��+j�h��e�������L�<@�k�����.��2R��j6���W��*nS?@H��;"EC2�+:p8���W�;�H���m^��;�}�K����B�� J���BdI�JN�@�K�[̔��s}y%�HSJ��v�qfA�r*f3�lx;���0mT����wؖ��xâ���ǨjK]����E[�j��ϯ,`�^ug���5+�]�ԻFO�Epj�>Q�������Df�,�����P���hخV
h,w���S�7@�S�p�n�3�E���hb4�Ke�����-�=0���KO�b�պ9�Y82�E%F��0��Q��Kgݎͪ��־�$���e�+Ø�o�
Ǫ���!$ii�f�n�W�`]Q��}�O+li��Z�ژҹ���쌎�V��];�^�X������Lv�%N~��hM��HCm���w�����M:ʈ ",ڴH1���ޭ�s���N��R7�=���Ea9j��a�~���-r�mL	[~���6�f`�~��EKU�OZ^Jݸ a��.�S�������8��ԧ��ֺ&n.j��/[�+��:�⾪j��-�{Ξ���JI��@pX�SE8*��"�A�*���d�_s�EIZ��u[���^`�Q��V6H�|~T�ؠ*Rx�����bHP"��������3���U��;�E���JA*J������K�閠3�����j�]�~Q�}N湁^	��S�7]�L��.w�t"#��Y�h� �Ȫ���.�߅�͞��aW��D���?�1�A�W����%�6TS�+� ��b���d�I ��p���	W9P�P���U�U��ʐ�ӌ�[��x���M�O�##�D��бu*]za.�l���g�/|��&�6�B��M�����B��P����#�y�����W>���SXZb)p�Ԭ�kJM��xZkLwQ��d��V�U\�L܀*ѭ��A�VVq.CaM`!y�&��΋����2s��/v�̻{�Ly��Qxq��b�}��䲦L)����
�떍o/���}���6�}��$��(���E�����^8���B�c�/�/v_�����j`�\R�r+{SD��n�O�~�\�5������:^��*@SS�#���8���be�Υ��Ũ�1�6�	��hi�fl���T�N��AV*�����6ˉ;6y��43�A�$�)�j$��������H��8�Z��$S�lh����%�uǘ�qE�l��E��B��uY�0BW�E���kv���S$k�����^>��\���s�A7������~��w�/H� �xc��$NT�f�r�"�I��;�W�<'�~�;�,�ܜ	�^R�@�P}a�2���54��D�B>WX����Y�lF���}a@��;6 �� ��qG"�ֹӺ�,�;(���nP���=��Ӱ\�/�W��P%^�$��1�$D��mh��p����ۊ5a���~&�&�x�-�fNn�c�����C�'�Oم���i��`�0Jyi��B��
�Q���y��6�5�8I{�Pfo���aq��?�N���m�vc�-oER�pU���'�r��g�Kh�t�����'���zd�2�P7� ݺ��HL]V���X,�on��̲��upQ��!3�	l#�6,�����B�//���5W�	�.AB�l4b��f��#o��oLxq��Js���8��i�W`����W�X�S�d��G���u+���U���s�e��gZ0��3����O��cݭ�'���Uî�ڰCYW��<[��o�$?q��l��>P�t}� �+gs1s{E�xDО��|��K�Hp�!fYk �_�ͭ�j�O��_�7e��b[��4�����J%����M�"�����P�8�<tv`F��2Nc;Vj{PGK�p"��F��:��0�����>�O�*��v�䤺7�`�tި�ȑ��:�m�s?�H�p�`��K`��n}�Q@�[*��@�g� 骩M؟���_M?}nb�
F=5���eE��u��w�[[sۈYn�S}��Lg��D��t���/=ɲ3^+^Ha�K;��=z�އЧ���B<��U��2��u��*$"+����z��7JF���O����e\,�S0�:���M�K�G�n�ż �.�%�w˱�u�Z5�6��Y�D��Cov6��ַ�� K��s2���N��,����p@��R�zrh|6G�\?sd�|~�pc��.u�(<�s6�bD)k��E4��48f��p���H�B�@.�j�3|Y���Ý���ib�%�-_B*RnK%�Y�N	V�[}Ѥ�����OW�>��O�������s�p��ڊ¢\��t��/��D�L]������1n�v��;�TfL;äZHݏ���\5��^eebn���h����bgd��"�d4����H��+ќ�\ �-:C����딤MEP�`�I�"S�76? ��ZnV�q�!���F�v����bDb�DsN�)���?��;O=��gc���b�&<ӁZC� V��&����2o�VT}<�,{J��$�TJǰ�����<���"�4�]��r�m6��� �4��~\����
�z�:qzr6P�X'�����lc� ��h�d&r��렛�Zt���.�w�]@�$/�(q���l�����Q� �EU�p�.մ��H�^v�\�:����w����o��5%Z�P�Y��`�� 1]�i�xҽ��gT���4�Ҕ���B����5P}˅%��f�����6�*6��OX�����>k�̼%+�^��/�{�������F�X��VE���L�=�r��Zd �s<+-֒���$�
�!�T����0Y��5��*� �l1۔C������+�d��ͻa6��]�[�@�_�kW�9�ɫ.@��,Qj�����ތ���zk"�^ф�t+1�U��4z'^��H6*p-[ ��gi��b���::ƌ�Q�[s;�G*&�Υ�8�r�����4Q��$�gט��՘�Cs��ð��p>��y�JI1�G
[瑁��n�����K��Bo�˜	��T�2��ay�*I3�1�0��.��M�=�w���qS,��)5]���$?;S������hcx���o��(]�<S�H���UÂ���r��`	�G����nd�g �{���	�6�KO@Չ�����n!�$�Cؾ�m[H��Gk�� ؜?\���0��2���x���0�8�#`b�L�_'�:�+;���A7�p6������e7~vڀa�I|y��j�Ž�a�8�u �Y#=�z��2��Lr�
m�]���]W��F���T1Az?
�RK��-F�I���v��7T�����BӅ\#�T�J���4��V6�MG�I�
�(ҫ,7o���n��4O?+RKʘ�F���<��(֡Gb���_���Â����<L�){fWX6��5a`��C�ٺ���^hV,�����r#� _j5C�Ƴ�,���eV� 3�y�)ߑƕ��F���uP���~;C�\r>�����u�����6�co*8[]9�t�֊�����-\�q���<�Ip�.雗��F6%^�����y�$A���B��}���is�#!�ea5���go��Ў���#�l�lf���KL�'3�7�~u�n������a�G���|�ܑ�j�p��(u�����O*�;�����4c?���*�%51c��n�\�@9Q{]�z
t��vM�#X#~$�a��/v����?���u&�������,#v��K=�c��3��� g�6�c�,�&T�mǄ��v<��jmW5q��칯 ���/,;'��B5�[L0���ˋ�U��;tI�j#��v�.�e�`8�}m/��]���5z~}9>Zz�l�E�*9'���E�[P|_���B�db	�S�.�{bܠ?�a���#��.�䧩J���/9׍7׌-l�����!�K�(-�rC	yu����e��C7�̣�A�����(`�̵�8���|)���p�C�\X(�I�s�M�D�v���{-�\���E?��~�A�!��w�dy�B��e*��1FM�����20����d�|�P�*-��1�\^�Pה�2�Et�G���Eb�������5�r#�58c�Dc�c@��v�좾	kK��Ϊ������0�g��gs�����<��lb�s�u�=�5$��^2�Q������y�-J��WQ'-���w]��]|�y�k�<�@��ʃh3�~#p.g"F��h��1� @����`�f����)��8� ���i��˸�%���<��� J�eo0]
)TY�Z�D<V�ڊ��zV�&\��#�cѱ\O�q���H)c�T�`}
Qn'A�Gsԗ!�$����*��
�ƗH$0�!=c�4}gIW  ���	��U��`��j1�ի~07�c�S�K�� ?�_F���J=Uh;��iZ�_�T����U���ޫV�м�.��0>��;���ɛ-BM�(�{�_-y
����I؇x�iF¡�s�7��A�B�WE1�y��{8�8ly���K��,�����EFUN�_�m�I�4��̍:V6L�����}d�n����+=�R�O7����FAO�d�u�����k�r�F%�����g�n�ʫ�cy��sMڳ�x� ����K��\3�c�/Wަ���T��~'�Qi�Z(�VYNo�?�O�R��^	��V=��������^����]J��ƴ�U��Y����m{Z�,jXށ��<T4��"ʑ�u������P6���3`�K�[��1��'����C���M@u��8��[��Q���_�2ϫ����b|��oD��~��/_�|��W���&W2�nhb��@�+� _b�GQ@ye�O>3�$v9�822� �T0�2� ZѲ9��H��֊k� i>�J�*
��9���D��9=�6�E�fI�7��R�-��u�1�
�N; ���)%��W$q������З�Jn�A4�o���J."�MG+�߳���p���~����=��b˂�b��a�j���˧qBMݘt[հWFWJ��j�L\�ۙ��]����^���/�=R��	M�*$���G3Z�M�-���^� ���¶�=�����[W��W��G}3�`NL�p,vH����c:T+���7��hѩ?*t�ʜE�C��m��"M�$����>pg/�q�(����ڠ�]:��37�gy|�q�Kժ:(�9��KrX{�	r�
T8��bG�\��j擻CJ���m�KyQ�,yL��,t�?{ڄ���zYI��{J1����΢x�F��L��0�iYQq�X��;A|{�M�?���0�D���m��C�il�D�d�.�����X��8r,�u�Y��%�w�g6Ei���`�*�Ł!�va0Y�wPr{Ň`�Z�}Ӣ.�����2�(?�Ĵ�f*�qܝlA�6n�4�v5�FI��ݖ
��k̳Ƭf&=�$'�-��o�q5��w"�o��<�l��S����2��K��+l��F1kEK���*s��
�5?��_� � w?�B�`�A�Bv�t��&��d�%!C#�&k�����-WE{�/�b�z�i���8������+�B��zL�`�4��0g��6�Zq,pg+��=�d0i/��0���}��g`�y���	��U���GkI�<-=�Gj��y�dc��.���$%�{wɼP�h�dT���zf���3��}���p�}6�W�$7���	kX���/Jwы�ǜ��i,D�J%�C4gc�d"��+�̏�Dt)��i�<�&K�0�Hh���]�Rk#�1}���v^��wH��g>L2n��OP�̃$��L�v��3��*��P�dg�x[˗�⍦*�-yasp��	���\(
'�d��	ј�NI1`/H��.Dz8-� QB�jp�?�\�R�ĸt���)��������~���x-��\q���L��6���@�u4�����k���u��x��"��M��4zg0����v�t���{�U� �C"g�~�O�pY��8Sq��N����]4�W� ��&_PW�0j/���0�A��(vё��2�F8ay��FX��5��&��)@�ӍҌ�c=�����Y���� �Ū��]�ۯLro� �Q�=taӿL�Q���U�l�i#�*�9D�ߺ���J����uS�z�'v��у�]P�&��M�֞��Y���S����d�*�M(������|:$�y"�Kna&QLs�+�m�G�(WtH��&\X�L�F&��~;�C�H�X@L��N���Ȑ?I������ԛ�V.��������p�P�8�8qd���C�Շ�������V�xG��Q�Z��*(��|ٶRjmh+=�{�������F�����Oo��F����3x���/$��OU�?�J��]V�R�m9"������G�Ԓe%�v��a~/��?z���x};�:M���m�b����?Yş!�Ϗ��q�&G��KnN�;[�w��H�A���M�*��!�1�ޱ�s�i�E
��C���h���z�u��e���2祯�8⒐z쎿�g5l��D��U�7�m
����u�4&yV����/�,����>�ꃊ%�WI���Bdy�Zh��3�)3ܻ8���%K�x���7+����F�o=�J!��[���/��U*���嚬n'��ݡC�A'a�P���Wb�;hH1Q7�7燢����\@ޕ:ν���v�ު��ۆG�8�W��*�������h��.mߝ�Kw���#Z�T{k����������=9B�\�����#_��5�Չ3�Kv	�O/غ,�0����0S�gI#���L�������n	~�6��'��аpDX�#u�6�ԥؑ�Ŧ�K�a��~t�cM�jb��}��H���6�k�Ԇ�t!�\p�m�}wo:���<g͟L��y���[�4�g�-ߖ3i��l�9�:���+���<($L����j��M��<ki�Vb�2���j72�o�M�ax����7�0�74�C!liyPq����d��k�*!��*�.�x��[q<)�RUjhE0s��'x�D|Zh�p��E�/+Hk�BV�dXJ�9ƴ��ڷi�j\����21�
Z��T9����z�-�:�����&4�|��<������v�oMKyӥ�r�`-�k
7���|m�ܯ�V���ש��ܒH;����h\~��a�l�K٥t���^F�*ꟻ������D^:d6s��{f��H�)�7	exUK3��pb�^_��J�ʛG���xb!6�������f���օĿ��\�����yrJ��*��̿J��ɉ .bNk�##u62/�L��kl�iZz&U�ѓ\���dt@��I��@����w�����<��)o�R+p��>Escl|��8��h�d�dLN�Jݠ��aa�:�5���4��C�o��+��<�M�ڒ2��˄�eA\@p�Ne\�u�XL@/�Tep�Rq���􌊊����~Q���jv%ٞXp��I���Y݊���f׃<`b�҂G��.�a�Ԟ��i/�j2�+/�������9������Iȋ�f�1��#^պ�z:��u��L#1��(���1l����2���vͬ�%ѣB/�� Q��`_�u��=��M�����^K+����L��RD�4�௖�t���P�D��P>�t�g	8^R�,deb`���@�˪��J�$�j�J��cЈ bG�H�G�2J͊A1/d���bB��"K�~�k�{�C9��䩂v�&M^��H5�=� �s'@�>4��?�.����\I�2�8M_�>��=��2��M���	�-�H�+BW���.Y�����Vc�Tε�q����O����̚[ܘa�ܢ�T
�~O�� B����hح!�0<�z����m���΅�=L�:e�����+����Y���_B]a�� �fV� t֘��i�:H�e?"ri/YU�:H9Ɣ��u��h�1���7�ؙ��	g 0�ܭ+ ��5ԌO�Ƙ��ar��j3.�>��\/�a����x$�&ģ�w����fLR"���jX[�p$���IIok~���G"ٵ�O�a�+� f^~1^��Y��zҶ���
����[4�����M`�V����.�3�����2Ƭ�nE��%��T�>p�f��MH���I�Ʊ�'�U�gl�G�buE���Ү(��.��/���O��D}Vͤ����p�Glm�C��N����V�D'���Ã�W��:	��*K)�RG� ,�	�WE�9;x6&��}���Q冟����
m��gr�K�r��|N�[M���z9r>�⭤H���@Ʌ��3z�ɛ`��#�<���s`R;�-R�o����f��D���j�5g���9����� 4�*��4)�o�w��0^�5�[L޲V�HmC��Ǒ�*�E��<n�R��Mq��X�Ag��>�,�\��ԋy�j�X�P�"Y�u��h���٪v�3� HE{Ą���e��ݓ���ɨ\����Π�z������B��CV���u��R�r3Q��Q�sf̩|��u�	uױ��4/����hW��N�O�{>0  pU��\dϱQ��DYr4�}�m+N-E�Er�Lz�/�ӧ����Y/*U��%�MK<^�����?�%���g�]+�C�X�fٲ��$vi�"^���zy�BeD�r���x�n�����|{ő��2��������w��U���t��`x����JS�2�`�����(��M{=5��d-Ek����/�G�$p2ab)?�E+,��2�)z'R���q�<�E�k�6���S;yP�p[΃z�U `�>�su��8�����_�+��-+v��l>�-�I�ſ�v�P�ZI0#v���'�+*<зϰ��z�T�%��-M{�������D~����bt����ʗ%Z �_-&��t�𔡔}SM�ҁ� |�S����6:�N��\���Q����%U�P`�%���fq�IE�jj���J��T�>.6D�d�<��7�E͕Vjm=NȢI�[{Y����f	S�YfM�܁���XH�G���1N�z�����b�=��t�2�Z!�����"t��!���X�n�Xҗ��˛m�?�q0k'�m��3�l�O�'��-;�L'LRHc���P���kF1�6��+}�Je�M��x7�xc(S�i;�٢�.`�B������א�ss�PxaO9�m����) +�$����ٍ|���t⨄���P�!���2�k���J�0��n���Y�C������@���������y���	˨d{;
!`�DW��/P�!���Sv�Q�鞡��ǉ�3(�a�o$�YJ�,j��~���'���U����I��Mc*�Ƌ��Jh�O[��f���9$�`5Y=R���Ac�{a��� p�l�;7������ҿ���ٺ�8�P�&�`��5��?��S(�� ��f�cH��/Y��:�a0�O'��g/���<���`�ϲ�.������	znCo�!�$�(̩Iq�+�N�$�
��A� R�)\3K��.��#�T�84����I���K@.C!>�C���Џ`�'ƵQ4(jC��,��`a��(�Z�}-=�l�CyK�>߼�t�,]�Ko*q{��o�:�Z��d�tz�I�K5�D�7�]�Zd���1;�d%
;�6��� ��Ч}T�xٖ���(`_u��]��3�-k�Z��8�@��g�M�d�U%�[kMz���旇;��Sͦ�)�4��n�ч�bW�n�O��Ґ�$�g��?�l	���P�>�"@5!`g7�!Ę�T�[�c��6�G��
�֚J3��)U[�ß��yL�N� �Kvu��d)ʭ�I�����X1��A���t�_/K؊��꼧��w�%�����H|�q���F7���kۧ��#��# �ղn������i2�v���9�z�t��x7�~f���W�A�y��$���[�oh�zN=��������'�L��������FJ�E�x)~Di�_������rE̝{�	�����c����"Wٺ��)�.��r�o�`�|�O
;��Q���F���c��QFV��Q��x���)?U�)�l��fj�h��;���B�ۋE���=�q�3F��	���O-"m�3e���R�-U�TҷмoN+���u�UՁ:�[uȼO�ct/�4کnoX����n!L������Uk������~���}ڪvW��P��-|!��L���H�{V�4w���{��ETf�p�����P�7�m���r���z����ND1|̲ze%g#m�K���ڷ#Ч�"���:d[yrY���}Av�Mjn��]��Xr�_�Ƞ`�c��Z��%>Pb�h�48�X��Cp�����\�mkX�	��7L���§����H2^��D��C�\
ç��\�E�̺������#s����}�V�MRT�
��T�Bٛ�MM�Q��ch�ㆤ�g���TÖ�ӹ���b�F]r���!�������d� �d��$�@�<QPz��r�Is>?pc�qg�7���@�!y�;�+;�J�}.?ƥ��}=˟άX��/'�'�2&��|�VB��h����F�隗�33S��1aDi�/�����8��yn8 i(gr��?��Kl�a������:�΅@̙��r������tԺ��$����j�Y0Q�<��q��>瞮��\�ًd}��׋�����"��a��l�N�Zű��Iye��,=��ۃ�xp��ÖE8w����t�˞^��=����'��� 4I�`&(�A$+��V.�NfF����a��Oz�:���1%^.��Ҏg�`r��\�+a���oDU>�f���qP��<�
��36Y�x�ʃ�R�R�,`�������m��x���2�����̓@�[�u�Z01њ�i���b#8�:�V¾�W�����\ȈX��59��1��_��c�'�`쩈�Ч#q��`MdQ������LP�a(~���T�^��JgI��Um����V5�3�P����=L��XW>ևo2,^-ZS� P���Ę���丂8R3^&\@9uq�	C�d��}���Qh���֔$�*�jw=��y<���w�q�ɯɿ����PF~���h�ȶN��h�����S��x������L@<�^h���25t��
�R9�ECBf��{���I��1�-ݩ�jFs�G����ȸ�B�)��jgt<kRN��l|��L(@�U��O�2E�y��m�$x���nwP�{�6}�����p��<zҸ�ߨV��z�v�z�#�?���:	v9��-�c� ^5�z�E�u:~�"��ʋ��Ѿ�_i�.s3�<5���j�AФ�Yl	��a�x��?�r�q�Đi�h/����[����5�}����M�@N���2���O��[V�A��(�4+s$=!A:(N�#���*`�<<=�Eq����$��I��u�9�S䶾>: %�<]�(`tD3
މ���Jt����!��b%ʨw<��� 5����y=B+wfbaR(�n�0�I{��ģ�^% ���v9��@��+X�d�G�{4ˎ۳�ξ����!O)լ��n��u����nf�Ⱦ�dL�$�d�i�v�Y�L׊�ua;�0a+�*gӛ�]W����$DQXa��&f�zHav���{�x\-��]vF�3�r�~����+����Y�@݊�{�dy��W~�%�3��!��;R�i�q�e�����of?��E��햛A����5���-��0�z#�����Jh�W���A��y����4�F�y�ޤ��ֳZ�N��ќ/���gq-N�9έ�O�e��c�|�rBԆ����y�uZ".���C�D�/E�Z�[����]�u|�͗��n���)Z#�'�O���t,�����h;X����}ov�@��
z�{�~� +�d���ڜi��1l.rĝW� �jy�Y3���^: z�q� ���6
��++��B���Q�%�*ן���4,�����4m��&��X�1׷�w�t�vx#'G
jל[B�V�r00����r�/ �{0G���8�����9����H���y��g	DHN�-�9���x�͏�B�^i�Y�e�l��sWY�z����6\����V.�ʊhf귝
U.=�N�%y�Y����#���*�	|Q�'8.41�3�D�}��[mE|g�X�s�@�e]&V�L�/IE��V�u.m����۸ᐙ�gC2��^w��,�5��
��Cc��
���&l��z�Ze��G�/}1��|�`b��$*a��
�Q3)�����AE��X��
��%8$I軈׭��Ƶ�Ɲ�7�i�'�3?ǉZ���pB���o_=3S�&�e�N���9�^�����S�����V>y,�@|�n����0^��n�e��H�uc��('=K��������G�=�6n���O�D��U���A����<�n�E� U��q@�>/Ȩg���l)2i�`Ԇ�5�;"���9O���}��g�&����5(,F��dO֧�s�8�p��3���13�<��,��t�ﴥ�G����p8R-z������[բ���� s���5bY�O=��Fҩ|X�2�~R:��	z.Y�J�j~���n}�\fÊ��l�t,�T3�_���Q�����X"���߇���E�;�����g�-�~$0�W�=�Z�<�i��ٮ�@������y��ߑuOӣ[)��HR7�\���/���pft��Z�C������}k��t6\�P��Զ��u�]�Ω�n`Xb|�%�9SH"B}�e������2f�\`��}�
+.�����D`����O��o��zZs1|�:M��ߓ�2��hB�A@0P$k�H�|^�:|��IҫP��~�b�HU�f����3����Z�AH��qYeu���:���Y�g��{��y�O,
�� �Bؘh4�Q���d�
iZv ���ݮݘ ZYEA��6�s.���K�k�AM��F�6�CW���x�$�n\VСt��vG�Bl�h�r��(9:�Q��.])��4,*8�A+42*�r�6x�#x�*7�r	+%�j'I��oHDi�w�a���+���eh#��>'|� �)7l|�؀������ĞV�1��(u_%�p�US��6
Ւ��GL��l�|�F
�ߢ���J\��t�G���)�\ �/���d5;,���e�eտKDR�w��ᘷ���Ϛ������V�U$��^���Z_�堭a�y�i̺�IL@�N�e��D�q�5g�?.�I���?H݋b �#"N�%�y�q4��f��k�,KDq�����k�����	\`^�#�3`���i1�׎PD��d�^���F��d�n�
G�EH�Dj��sg����;�&� ��� N,#��yOQ�ڭ{O�.���')W�)�Uc�W�Ʊ�9��Y���t���v���2�D����G��@x!r�h��sڎL�>Z}���b�A��A��)�pZv#nvН\w9�r%���?�T����]��4Ar�� |�gk���Nn���&~@�4t|���A�Q�Ľ\%���e��I�w=�N�8ر���͙��
�	Ŏ�R;ljL}B"��Ȑ��"�.e���{���sD����BJ�O���ɔ(�<�v;!�������(W^�%�R�+���)E<s(ѧ��%�ME/D��y�A���Ե�uP���#bŋ��ҨS Ŧ��O��!�;���Y�8i�>�v�@�򐝒h�%�,��/�҄�;R����z,����ȩ�? �GvE��d���/(�f}�K)Ð֨J�;KE��>�����	ڽ_��<���PֵB�h�u�[�4�})�xjmw(�� �@v�(t����?� T(Mc<m��a:�E������O:�����HtѶ��AÌYB�A�TDx��vQ�������u�*�ȝ�I�_`�-+|&*9�	��ѷ�vsŨ��"�~n��9��\��Ƒ�������\*�c���d���W	9��4���V���ݓ�DLb��Nx�"��̯ur̄����K S���a�~�k��aل���1�ly\�Cx��w1!o!�6 ڷ/Y��i{~E�8i���Y��Rc:%T���}�u(�@�@�pR�<�}��}�Y�b�������w������|qBpP����_�)\�PDj�o��d�T4?�ձ#h�:3����PV훛U������[7���(�fy�(�"��@��z��hd������~��U�.�����#}M0Mt�.�88�9{F�DӠz2����]^�J�yc��Eҹov��s�h�]W�:̈?Ēc�
$W�0N�f�F�(-��������O�|#}� �E!�z3��Y!<��j�<-Ҍs�h�Z��iN`;y0jw±-~d�(Y2�K�9�� f�[D�	,�~�n���<�Zjt
����ܟ�l�6z,�t[��?�'�6�z��ˎJz��^5�M4��3���"�Q��(NH�]u#��+^�#Z.ө��>�l��O�j�y���,V���@������;���[-/*�=/q�|Kw�w�a��=Y�-�2]b`H�t�&iʹ�?�#��j)΁[rk��R�nn���%�2�*�����f#B �X��%q�s���N��|��ќ̭͉��2"Ժ�q�"�����#=x+�~��x7�{����(�hwSkd��6;0�����Δ���;yq�r���>��KY�8�%O<����d�Y���
�T�a!*��-p~�oHL�#�۠�Im�:��I�!�!}�Y?N�V������'o��_U�@��Q��Fw���o��nәDN'7T�u�kAWv`�	�YJ�VQ X!�g��
U�Tͩ\�c��4T��/*�Ge�;+l/�%�C��z@���ĥ�pՀDYrk"i|�"��E�j �������-�>�b��$���{�HV��4�5��b��a�Fϊg޸��%�iB24��k6�!���nI��&B��D�Q�)(V~�����k��u�Ǥ�����ɣ�z帺�G�h/��`�=C�S���M�0�+�Ճ&�9�#�m�j_�㗯�l��-��Ά3a?��� [�F�s���˙$a����j��p4�r���7�j��g��jjcV76,c٭�Ԭ�S�޼ʏ�ͣK�,�ܒUd.�a���:bQy��o�7Ǽ �+���D�ߠB���%����oqN��?̪e��^Z��k(���x���e)�5H��i�b�)w+��%���w�Jyc�\ܞ�*ל�:�6�jw���ѐ$�R���X�Im����S�cU�L����Rr���8�vmh�]��s�X�5i�>/C �+���4��3<L�|ˏ���&�6V�0MucCE�ϑ�z�LQ�sO��"��_�p
ǧ��A2�H�DL+��������e���/�L�/S������4�koUA �-R��+j�S�<U� O���5�/I���ST�uR��#��g�;3D1%I[5=#�BQ'�T[3�.tw��!a��(��P�����=�
�EXZ��n�:�؀*���-Cl9k*�L��@�����$ą*�Π��I��J�;��i{}�8$�t���J��u]% ׋N'�-?HuAIpA�{������I�ͻ�`:-��"�)�ˮ��c��z�Ǩ����PL<��vYd568������D(�@E�7 g�G�H�ph�< ��D��	�º��շx���$�dK����Ѽ��r'�h����Z�u,_���Π���^�>f��;<��z��tY�}�2�i��p��=dOF&�q���7m�TN#�ږ\��+9�r�T�W9H������C:�Z�{�W���E��qX�$��I�������P��l�X��)�+�x��<��t}Q6�p'��S� JyE:��c%���*J��T��ԭ.1^�j�CUO>0;-�֭Ĩ��n�oɷ�j"�5z����?{��6�8�(�]TyD5{��0���m}����Oj׼X��毴����ꫣpK]@��,!	Y��mó���:��$��V��l��<2�W��P+�{IKH�;��R��v��=)Qw�HH��J��I�64@Ȱ��I��*�t1�t�[w-�$���Dt��$���\C�yP+��� �M!9f��
Ϙ�ą��z����+*R�I�?j�������^��,��X���J-�=��"vMJ=�햇���O�1,��b��w.��"�U�d��oe��&4	l�`x�z�P�n_�m�W�p�X��
)Xr�:�8�7N���B�OƷ�n�)�[�A2p�a#�DVg��@8O���ܚZ�|%�A��\J�M�#�^' v!�/�-��o}7?5���P���Kz �F,G�[�ެ뷰�_�I����������`2��0�H�}��"(�����,��AŅ>9����U�P�3k=q�Db�{��=�#y�
9���"|JK�=�|���g@�U(�����ݖ�d{��%��`t��K p8�_�����f`��A�Sg-oqvWr�.ɜ�^Z�-��J�D� W���+��d��EG;�������	^�>�UN�6�%
�4M�߂0�YأY��R��ѥ'�E"������,ܪ�,n�5��E�P�>���+tM��7o��5r
�x��G��\+MU03a����!�qy���q]��T����K,���F�PN�K|�O�1�����sSr���߼��T�>k�mr"1�|��m�Uf)���O�E7�o��������E�3�P�/�1� hv��<0>D�]��
(;h.�,c��X�%r\���o����{��r��$�J��S��!�],�v��=
UQ�B�p�1":�B컱=-?��e�h�H�%�a���7��U�O&���\�z=
�,�\�}��8�g�M�t'ݺ:ΰ�Ë�X�b�(7�%�P��KŹ�j.����cuUu��V�qw0�x��<Y�'�aN��.��E�P���@@Cl�?"?�l��HX0��O��[�z����J��#�m�Dw�V���~�+H����֫�����|�oHT���x�i��W�B��b���_6�.�����w����Z�܎�tJ���U�㏩��10���E�i�ժ���F��uEQQG�����pL�;��g���z~�7�	��^���T��7ODIi(°�ڳi�"|�vR��mQ�F<��9�����ВI8[��a�ٛ�P��s�ɐ[(w�i�F|j �8i�^��yb��1�NC�ѻʵ 
y$�\+r#in����uِ��;@^)�݇������q�(�
e$Auf�-�>�N��D����q�BD^�	�Ӧux��E�h�Vd�CM�%+��1J�-*!��4S5��,Gv��䅭�
�:�z69.�M���.x[�f8p�gk�h&����&»������ϖ��z��`q�i�q~Q�=�s���2$�<TΚ�q&�Q�\�.H͌jm
.P{�3\FJN�t��N2<n������Ʊnw��]"|�B�S��@�C-,�٩)��hĜ�@�k�	�Wn��g���$*e�L�\�>Ѹ�H���@�&�O}�*�<:��(���L�YX�4�R����uݧ�J�,%��q���܁��B�a��v�9���gUI������K+#a��[\��ɫ����Lq��}��4c��%�w*p*�=5Ʋ�{e�ޓ��h���2�}����k �[4!��%{(�Ҁ��gۊ$3B���J ̖3�灻�N�f���ԝl�W�1{�Γ,��2!���s������������Ҡ80<$m��(�g �R?6%�p8�c��7ʋ���_>���++�~�K2l^�����-T���2���l ��{����W�q���É�K�9����4�Hڠ̑mD�g%9���4rD;��X��T^,���,�}�i*[�z9�I�*ƀ��%\|�ʯ�;YCޓf���4Ε�����(�c���&ϫ��&�o�ml�"�!;]ڀi�rgȧv)m�������\�.�w�,��Eoӟ���8D�gn8��"�j�i��lS��o;b��[q��F�Oit��B��[�<�ĺ��P�t�"���I�U�Ek��'�(Kc2n�����R���)$r�����~!���47�������M�2:���O9I:�Ix(���)}��\Ee��M}�Ƚ��25@����A]%�Y�
���	u��0�,A�.��)����-SH-=^�a�v7\-K0/��1�hˇz�FD�	�|>;���������%��\`����ט��[J^�yb^�g����z^y�L,���[�_q�q�ٌ9�����(���'��j����m����ꕦ �rـ�{�4̇�Mz���vY��~����x���:�k0�*�^���?kN��u�>�eX�4ԃU�K1�����&�ʳ�̻�e�}���ψ`T�Ho�gǘ����{C��fhu���pp��{�{�Ƞ�LoyZt&/q܌��0�����H��b� �o��;͹�B����qn�"ܿeS�ч$���ٙ�%�<T�bmW\�HS��)���3���=P_�z��`%�a� �U�sڠ�M��:_�՞ذ,2�����XԳ����K�b�;h��	�}v�>�CI��A��HX.>��}�R��xo$歵vC>#h/l啙�~Vő��iz5,� �����FM^�Eb�=z��b&��,���N*�y��L����]'�Ge� 3yq�@q�ʲ���p��S��)�`�R���$7G�Ā��^�7�#���Ȍj%ޑm˕��`�N�v�P[ƠHR�����z5D�5y�B@\�f�'���E?�'��2"�{�e��efZ�F=�����l�:Mi��7���b�7���&E��#��q�@�/�ƣ�_�8������VW�;y��&\�v
/\䭞�s���ѐ=�a�.*�X��a�p�%�JP�f��Y��3Gu
 z.2W��/�ս�i�������t�s"�:
�+��>sτx�y���{��Վ�"⡁k�~,�>M��I�r#�����Y�T��#�X��/�d��jpGb� �[�Bp .�.p�ARhI��͛���N��&�e�v�}څ?�;��VƗ���;�l&"���Pfv�
ET�o{,u��=4�Uc��|	ڜ�z�!Q����BP ���D��׉����)��SŻ�	�ހ/`v\�+��u�
�nr�wry��$J}�h�*�]H�؃����*�J�6�ED���,����)����D�^m��zP(�8�� �r#���1o�MS��Hp_ �U��_����[��+�gxߌ��߷�M�,�f��QD��C���`��̙@r��T#�f�t�7�`��`觽��,}Wϡ�v�n~���z��ͩz��Z��k}Uc�U"Ul,���0e,��d����ѭD"�M���t&V���5��%$	�نpF-& �'x#�)!	���G����"b�h+T�\砥�3w{��p�;����1�OAʄ�f�ѽ��?��)u���6B��~���EV�ƏP���=}�8 ���	�pB�Ac�"~a����l(WĬ�N>�#�ƌJ�l��̘&u���!�z��"hg$�͔��*KԜ|�b�l�l�:��y�=Q:z'�?�?-�mܔ�E=e�'�h9X�r L񓫟㎷$��9���v� �d�`�%Hw}�Re�!�}XZp���˚�����"�
E���"��1d�� �g�`�uO��I��/�|	� ��x�S��etK�B=�6�yxKo��+�:�:�Y�[�UH��+"�n�;��W|��|�׍�$��/�IتE����H6e��*q"�K�kN��'��1��Z"��6(	W�1�rI��MNӤ�TQJ9�l�����r�粓�B���A�iꀿA�-Θw~�`7��͎�ӕ�72D�z�$�L��X�jY!�#/��b(����$�X�b��ZGn���?���a塋!�k���Q:�(-H
����q�n� �?�&�5�fy�����ds������o�Y���}ܼ@[����))(��}+�!�(G�w�l���VW�f�3Gd�h8ĕ���V�m/
X�\�<��䊥�j�����4"	'�楜aF.�^��7����Q�ǃ���Ngif��E�ERMy�W)����,�����H�����|��1tM��j\x�![1�r�\�4��~�7�/V�sg$���4O�hׄ�Q���`m�)b�/�zL
J2Hy(;��V�a� і���(��{����n�-�#J.*��iVk�O�B������EVJ�!��ۛ�ͤ7�YF����=x���w�^U� l�#���5�����A��eD� K�����-�:(-�\��!�5S�9%"��+�K�+ӎ�o��������Ҷb���@j'.�b���]�c�[%U�G��9���佪$�UfD}��͵߰�q���Ț4ԭϙꭆ��6���-����kJ���*^F��S�H�[*��Y��[�WO?�f���^e�wA+�o���4�����j�I=� �i��M�!(�i4�MU�TA�vP�KO־4�����᛺����g�,�����j���@�*���k���E��n�	�����ש�z9bP̨@]�����h�k�Wa���&d�����P�n�#G�{0 e�r=�\�s��*P��_�I������u�<�őV��W�r��{8��D��w�>�����b�y:�b��,�	dz5o�'�l�4�b
S�L���]�	�a�8����(�
�i29<JY�k噌��t�ʊ��,z�Y?&S�a)>t�=�!�](>�
����tNY�\�^�b�-�e��Q�8�W��i�'���.#A�U�r0e�?����v�\�����6b8e�Z�����#Ň��K��T����6�lº�z���iC'ϫ١υV�����$H���H������WG�9O�<c�oS=��"Yq'��1��s:�Shf�p����Q
�o�Q�����Z*���v@;�O0����Șh� U\B��Z��t����L�����Ek��K���A �l�����w~
��s@��-k�p�5F"rD�FS�YX����IXif�9�V�0\�(C��} ڐ���M��?1	%��污�=���;}*Ƒ�\t<!�4�d����8[��˶2�Zvy����~��o���#)�;펊��jN���G�{��2w���๴v�r�m��l@�KiH���`��T�_I��_ؾ��#}�y��y���$xե�0!�7�Ut�j�{���	��z��:���<���[�����������l��Rȕ��[R�+gv2�E�jw��)!�.Y�������վ���'�8�&+O=�j'���]��B���/���?�u�g���]����3	�ca`j�#�|;�����ĺ�1�==��gk	���l�F'�ֱ�"C�E�zS߂�5��ض�Gx�2�%��=WK.g�w� ђ�G�e`U%4��%~QW�S�H��ed���b$\�!���,�$M)�i�l	���cJ�n2��w��b������,N�)w�Tи��,�v��=�_$��b��Lhv�Е�va�~eZ�w,�JӺ����IA������i��}�谼�*�2y�4d�k��ZUwѯ���S�v	���b��1 Usһ,�r���B���٭SI�Gуa�LS0w*[UKL�}e��u�g�$�4G�)�t��=ux�J�.;@�Ӈ37�F.����3W�{�$�һ�S�#�1�\Z�R�&�>��r2��b����W0�:ʉ��'�=���T�p����#��(fSw�����#�x\��O�����|�W%S��!����W���jg�ϛh�8b�U����p�csQ�a�.&Sñ�T�Ƨ�8�~����!ɹ�e�f���x4ʸ�te�Eqoʥga���G�H%�E6����e�3A�k����A���-�'O񒁎�,B�d�����O�ݖ�E����O�ξ�tBt l�Q���m�q�v�N�2��Ў7U����:��7uR�����/�*B����[nRy����jĕ���Ց�a��컙�֌�5�h�+�Y��\iC��S�=� �T)��&��r=?��E�q�&PC#/�[�0�ǫAұ�a�o��ZE�������3=@p��?�]a��AP�D�5��6���}�oU�E�`ԛ+����Z��:�IS)"��f�5�4�q���_p��@�)V�6Y.���8�`�,}=ј-�o�I��1����`����l��9x$����]*k9G��R�w���������ze��	.�����=�_�ҴpM{y�����ؚ9���~T$H�2K�؏Q+9Pl�τauJudt�&T)�h��\\h� Ltd���1aDl�a���b�q[�8��zkFZ��R?��mI��q��˃|.����t���ޛ����7g�;Н�U��:C�f�t��D�9�M��yP�پ�������(����'<ҙ=�P�qmR������s_�u�э�OZ�]�s��RT9�L�c?
v��N�{&r2t�WdұD�<ѓ�j�7Ԯ�=���ʗ���X4�b��F���ms0�S���Y荕l��	fڒXv��g��1��t`~SUJ7�]y��!��� ����1K�V'R�������_�=���B�g|�|��]�V�ϸ��u�58��1�DM&9Y���ƪuح��z4�u�<)Q/6���M.$t�#��͈|���Ƕ���C�w��jn2lD���:�?A��z�@$�P�L8[=(����49����r�Q�'��XZ\�DFqI.�\ �=&�9�
��a7�1��x<�O����_����s���v&<bW(Q��}���D;�����y}1��b`��Y2�r�+�.]n���WN53��_�Q�[.�>Y�/ui�pφ��V�΀�8��,S��{E��+�;�l�����<$�c�`�b�l�Ƭ Φ	9���?������B��c~�1&��$����F� �"����rU���d�7* ǀT��-A�xe��Q����@�������ƞ�-(}�
=o����#:��<twm��d"��F�ӟc%��QA1H�ӊ4��sXz����(C�:�kw�'?TǮQ9��Ba_E��h-e!t(�Xt��+�_�>�BY$?�!���\u�0�������v}��ED�7s�#&m������(��D���x-�ʐ
���܃C��2��
�u��m�H���k���T�V蠲X�S��D9ອ�H9�I�Ğ&���1.\��C�䘏�?�:T�߿��[�|é�}���΢3A� )��p��ˈ����~�R/��7�R�V��c7��u@���
jf�[�k�(CF���� �����Rzo�c�XM ��^�@��3������ѷ�87�������Y@��O!�Db��]���e���*���ǧ�<G����v@�U[A<�6��a0����"0'�^�#�9��^����Z�{p�G?��sT�����}�zn��A������R��_Gͻ�H�� 4��l�F���<�}s���'"i��>�1P1ob,fA��ʛa�:���I��n�#㘮k�x.j�Ah���\$�~p�/�YgO�l��z�ԅ��qN����m�\��S����[�\��X�����Y�M���`o��m;x�R��d�4�ܕ��|^��0��v��.��iפ����>ΤB��/�[��ȋm�2=z��@.�#����t�xl4b%ɢId���yL�D���g�+
w���ѽ��.�A���p"�M�zĒ���e���JJ�[��FQ!6�uʍ�*������.�N���r��c��&#�u�wx8�V
p���A�����Ԫ�E����;T��
�k�����ӸT���YN�����y���!EL#={�� n��ߔ�a~���z��l�u�Vkd��-��� p���������f��E�)��Z��yeF���h��)�V���8&(����W�a�Z����J�;�	��v�`�ړ�S|S�ӓثO2uc1�!ETs�GQ�	�cw��4Ϲ�֘����OdB� #i�|B*A4�|Yb"߸Z�� ���r�&O�����s���J�¯��~�%*��^ʏj�ZS��V�Ib;D�0���ų�: T�������e̆�Y=�j�\Q�-Au�k1�-��q�)]r��}��ǿ��)�X�r�ߎ��
���,bױ�2����<!��T�����g���ȣ�ѐnQ^vu;yg��b��Y�r�����u�v�[�rʶ��/n�+�k�V���$���η���������[W��W�'@�:�:��LG���7}��������M��z�U*�UԤ_k>(�8���5V�@��;����п����M���uMl��ܯďX�#��"�L'H�-Z�9�"%��\�S���W005��V˶�8͑��.�@0��#N���	�� �����*Ơ�!���
K�����I@�r�f�]�?i�rሤ#WZ?w��o�y��58zٝ��j�zr7Yݵ�Р	5~���ҝNyk�)���R��n�5��Zgu�ܚ��q7���Xj��Ll�j�)0�Q�'�H��q�tTx*Ô��9��t�z5��z(`���Y�G�[�F��f���E�����^��Ŷ*������*�x½P��U���x�
��e-��h�r�ϖ~��e�?>˼��3�����o�Q���=Z�_�-=����U,9fQ���M��iLI�`��M.D�	���א=��0y��]�x�(N��3R�,����*�u���^�����^S0�Z����tRa	:��*l�m=����N ��owI�{wm�G%����|s�b`Sz%��L;��$���1��	z��o��IHz]Oۤ��ҧ�]`���C�|��4�3-sS��j�*r�g��yB�\���.F/� �� �9[�� �N��q�,���c��&�֡�n<fn�:1�q�~p>��'Dڃ��~�fL���B�m c�~h��*h4��z��Ӡ-��i�+�S�r���'�~�Y�Th��>��x/�d;�Cy�9H�`�Åq�ط��.l]��u�x!q��4�Hh�0������;������@+(��v�����z!Q1�x~0���j|�|�N����pi�\�I���>�ı�i�2CB�ϣAV��Kf��3�k٨�ܚ-�c��|��~ܒ��P0��t�n��-�_�A���kh��i���^U0�v��