��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� rā�SZ )����C.��&0C]�-��[�3�-���+��պݣ�k�J�vo`�A�����f����u�X���v�=�а���]Q�Wۿ�߸�=_Q�X����j>��Zw�K��SvX��ƥ.���#�����Z�0���#7{��\S$��@1I�QX~TQ�E��db����۰� ���>0�%�9�j汈��}��1� ��2���h�G��SeY�a���	'<x�p��k�H`�H�j^y�0�s�78+���ֳ�`�R3dW��_��{p[�?$�s0��#�zS�_��bH
�c�p�IL7]� |����Q�� ��Rr���=��E즕2%�����`�^��l�q-�]�p��jf��Ӽ-f%H���ȳ�>��+���M�71��4_�) 3�46h�rb�J�W� k�h~K0�>P$�_n)���5�r�j��W�J&޴o��$>��6��ŀ�;A~<6P��K�~��f��*I
�Z��}`q���ApC��n���g���3��-�іrO�mF���,�$��@�BI�q�}��Ȥ֐����î�䂧��@������U���vU������ �T#K@f�㯁����|95<@���+�-�)�����K���FI�k���*@�m&���
���ma1[�2�u�I�\�U�yu���o�|��2����;�W�W�}P�K>%5�'�8���׫=����k��,�t�M�0�8]q3���N���GvZ�i�+ C�e
��Ќ�S�v<%���q��e_��
�k�夞��>ZO7E~��5k�TW Aod��eE���G���ɑ-'���?�G$����ќ����8ɸ+ 5ʗ���l�d��,�J�
�^�3b,�����J����#n�zK����z�&��;|�\�^���'e�W�����">�w*	FO�Δ��v���I�h���!qo1g�ej�1k���
b���P6����lIy����F�&
����4ps���#���o�$?o3
N�'����9k��X�h�����2�G�Oƞ�ۭ�6�0i=�~1�n������Y8�5=�j�� ����v)x������
Qz<�{�,��$����L�{1��wuڭ��Y��QVC
*\�tږz_Z��]�E��1$�b�b���6�04f��/x"D-�����9c�L�!tΪ�7�{��ݱi����c��܅7	��ʏ]��;w��-�љ4�կ�%�C�ݑ��wte�Ҋ�:�h�,_�����3Q���	��oǑ-����I���G�-�\%���B���_{������ uK���*42�H<ԁ��<#-9!k���)k����t"�X ||�5d^�(�'pL1rsK��)�$Ֆ�x$J6I��>�Q�ĵ��V.W�f��j������5G6M�뿹��'d�I�R���#�j�,�"��h��S�b���AI�Y���`���E��fǞD���'�6�~��(�u�.J�T�/��
�9���Uv+m�����Ü�aL�W0j�u9��(�\N��=S�ֳ����F�Wc����ޛ������¯8Ҋ�qD��ZN\��ao��M�M4���nG��P�6����L�=~q$C6>	<@qc���D�
�Gs�?��/l�rC���Mn��Gu��z"}��gm4 �Ǚ�X�x��#���rr�sw�1q =S�:0GB�Yk� (��_��}��>	Ư�<`>��|��J�`���U�i����+�ȣ��I�ּ;���,��{8N߀^�q�M��(�ixq��-��� t
��d>��!`�B�T�Q��.��Ѣ�BA�;{�ju�:/�=x2�5�l.$�(��U�j2��8b
�E۝���O�E��4��u�,��;�n��Q��ݜ�MI�)�Y������N���]��;�;����=g ���i><��>ɒ��L��<�S��e�F�g��%�  fh�����o��0��������m�co�lw������[�D�W��ybF����ɵ��PSYn��V������NeD6��4Q*>s�z��V��XQ
ك�ec>*�)���F�U��ȇ�i���\��5��3*Jڞ��P=
6`KcXf�B����nE��J����2H�߆����5�2%�JG��8���|LZ 甼�B�ډE��]a85z'��5B$��I�����R��i�fF���}�'R6��#' ��N��!��sJ��@vN8�����,ۋ ��k�81�����%6e=݈L�a�^9���i�WѦ�~�"����(�"�$)_����� ��H��{�BP�]��Td<��8j ��U�9��#��*�<�A�2d�j��q���q�ս��'PVxLn.9��/~^A$�we�'�����?X�~՘���"NG�Y���G�����.��q�œǙ�L9dB0���S����h3�%�<����N�Zlx�JՖ� H�C\����Ճ#�S�Uڽ�Q���1 ;en���I���HA~�{�TW�+�8ʊ'�QRC�������=W>f�)7�`�{ ���F�(��	�&Eb�f$%��+�"�$�r×/g8[I�f���+.�����\F&/tp��>�b������y=��bR��&�[�ϝ��7�+�D*�r-�Y�u~,|J_��;�iZ�(�AtO�gJ���f"���y�>h�U.2�-i�C*�#�'��J������Tr�6;𝓬K�� |j�9�??�7ںޖ��>�Vf����e���檟����u5O�\�����j�y���*l�JS3ax��bs�0Z�����=G׭A���O��q���2���%���I�A*�����A�0���-D@��%����gΖ��û!gZa��|_�H�+k!3胶���!���ؤ��1`+u��|���JK����R�-���+���1<J�y�>uú�0CǮ=�l��zߍ\	���\�q��i��±S���CM(� $��BX��������B##v�Ͷr�~���3+
c����)�M��-Y�5��A�炐]�	;���Z��m���[ ���T 83C�mRrA����(�nG�����nL�&F����G
�AJ��|M1�A%��~�\��S؆e���x��>���&~h�U�wOc]�8���o�p������:�ޙ��B8A�N�tT(��4u��/N����i;�ϬxOR���f���iG��ߡdi���^� }i��X �y�g^���m%`XP�A0�B �d`֯���Yw��N<3��4;1��L`�B`Vc?^g������~�(]��#iIwkk%��)��f�P*��د`�s&��bI�f�0D�v�`�����MƦ���P���ᦌ�����Hd�U�Mӯ����d�P�&vj�6р��#��Qiт�V�����ơkb�Ω�23*h##39}��8�A8��1� Z�db�(�z/JQ�!�_	J� ѽYs�t���k-�7�ޟ3�[V
��������[]�2,+]�^I�Z����0����	���-�~��e�rv SlnZS+ZF���%�̓T6�@H��Q�ίg��V.BpO@�P37�gq�N��j��#B���~��i�DP5�<����]WJ�"Z����r/�%�^F�E������5�ř"7!%���voq�R���W��t0u�>͢Ql�U҆w��/`9�B���9>�(	�H*�q�^?��zܟ���2v�*��CD���� �U��w�SaJ =;�����P��L%�AA���BXrMBY�L��qDB`M�������{��`'��h%�
�g6�kfT{�T�E�J�9�\�j�bN�T�h��Cb����^�k�����؄|q�~�pD���z�߯+Z�?�0rb�8��>���B�_��l�LQ�S�u�0;��_&���X
�M���`����S��n%�m�|�M*�!X�U�$<;�[@6�B!eL`�!oսô���84���������oY/�o�=����9Mc����!2a&�	�K���7b=�4�k9)��5h�4�;2A!u�p�mr�A%SƎi9�g�Ʊho4hZ���w�퓶ŷ��aA_�R_/k[����ǆ�a�E�W:�Lo�'�Ds����K{�ڻx�u��.i3D��2%>o��r3��ৢ�u[p�J_�F�d�O|��o�i>���i(�ۺ�3�}۠�� ���W;u�r
�ns�&�Ԃ&{A�I7��i�(hx��2��l�av4̮����?$(��A����x�����U
l�?� �T1����R�p��>@0������<�Q�kjy ��x�#�[#�5r�B&$KL��T���	N�P�QD�@�δ�/;��;|ހO�Zg�⏈~�=����i)�x�q䐟��n��=� �l��w�_`ݢ���'C5�ȄfG\TF��|�N���!������t�h"�:MI5�7�g�5�^��18�Ǘ���+���Gf�I�rLU��1�O�?���
��k�nI���R���xa�b Ae�y����~r[�h9