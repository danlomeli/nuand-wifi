��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� rā�SZ )����C.��&0C]�-��[�3�-���+��պݣ�k�J�vo`�A�����f����u�X���v�=�а���]Q�Wۿ�߸�=_Q�X����j>��Zw�K��SvX��ƥ.���#�����Z�0���#7{��\S$��@1I�QX~TQ�E��db����۰� ���>0�%�9�j汈��}��1� ��2���h�G��SeY�a���	'<x�p��k�H`�H�j^y�0�s�78+���ֳ�`�R3dW��_��{p[�?$�s0��#�zS�_��bH
�c�p�IL7]� |����Q�� ��Rr���=��E즕2%�����`�^��l�q-�]�p��jf��Ӽ-f%H���ȳ�>��+���M�71��4_�) 3�46h�rb�J�W� k�h~K0�>P$�_n)���5�r�j��W�J&޴o��$>��6��ŀ�;A~<6P��K�~��f��*I
�Z��}`q���ApC��n���g���3��-�іrO�mF���,�$��@�BI�q�}��Ȥ֐����î�䂧��@������U���vU������ �T#K@f�㯁����|95<@���+�-�)�����K���FI�k���*@�m&���
���ma1[�2�u�I�\�U�yu���o�|��2����;�W�W�}P�K>%5�'�8���׫=����k��,�t�M�0�8]q3���N���GvZ�i�+ C�e
��Ќ�S�v<%���q��e_��
�k�夞��>ZO7E~��5k�TW Aod��eE���G���ɑ-'���?�G$����ќ����8ɸ+ 5ʗ���l�d��,�J�
�^�3b,�����J����#n�zK����z�&��;|�\�^���'e�W�����">�w*	FO�Δ��v���I�h���/�*n
�}X�ƪHʀ��!�w���F��n�Q
����?�Z��
��	�6�ؾ�^q�M�`�(_�����+�Vd������k����ey���y�+��������ſӷ�c!�j��Y.a����ңfL�t"�3W��mQ<���4�J��0� m(WLt��@z��H#���e��V�Po�c��%$�&��E�u	:Q�}=k@>	P(�%��%劃Z���x�_���S��FJ%��b������x�J8�ж;3��w)�vZ��w��/��i�3�_�d|-����A1���b�	�ұ(��ʗ������X�������z�s�:�y�%t�2>��د%�z���S��&��13`&�~D�6��t��(#oܿ�y�#�����Ӣ������� ���������ʴ�G������y-im�D,U�#R@�0S�m.%�`k��aI-����j�)�1�=�^��!�mrll��Nl�4�j�̤�;1��+��i��"�	�t�k$��b�>iK�w�ӑ�j9����D�
LӺ*q���%��1XC��RS
I�t�m5n����;��=�1��`[����h�+������"�h�s]RD�d	�k�_�p�)����&}?�����C��_FEF���d���E|E�<6�)��h�B�y�{�l�Bp�T��$c�E_:�݊W?+7BrW}f��M��a��g,1�VN�����FE��(*s����p��H0$�^��"	���Nީ��Y�(:��{��er������h^���*��s����\�G�y�矪gЮ ��[S��2F�=�������ߗb�A��/��.��?v\����gM9q�I���q�A�ViʿD��ڙ�c4L�%�D��<'d�uB�aȟm��B/�.�+�x��w�|�r�`��+l��J�6��/-e��x���sj�R��e'ү�So�T��*��6x�Fy�s�J3�i�kZ���"�%�l�:$�0@A=c-6����t��veL��<��K%.��R��1�������"M�}V�� ��G`�6���(Ĭ�u3�������j�#�lŉ�jp�.��
�����{L��8Y�Py�8�	3�_g�������/C2�\���O�h�5��wc.㑊�ٓ�a�HL�Y?��;�TكHҹ�/5��j��"Wv]X���h�}��$6�3MM���:�:��ڡt��9z#�P-'�L�;�{������n/���v5����]��@�≎����dta���W߽����|Ϩ$�<Ŵ���)77/����pp�t1?�]���A�P��*p�:�`�Ŝ7��͉�H�#���$X�|
Tu/������b �����o�й6��f�+��(cI�����v�����R�Ҷ�Q����J=-�}�'@�4)�⺲/������(�z��;;�7'��|b_��5�v�����03c�=���1�]bV����1h���uO�B��<`��b�z���Wa�4��}v+�W�@�����&�ץ����jk�e�C&NA��u=)�r1�q+����n��1�-:�|�LU>�o�.��(F��#����|)��6��W�'�ϊ��4�z`2�,�C�'�	D��6!9]�����Y�T4����%�S]tNA_ո�Q���=���u}�f��`M0��]�J��l�Jw�Re�iK�ŵ:��V��\���Y��
쩧��je}|�S�:?�����jƕ@�P�3�����
���7�Rs0��G�^�^$h�DtI��<)�D�t�w�07���Cw�[d+���/0� �|�H/��ugc~��`(��o�v3���.>���v��f��R�`�/|@LFҶJEݽ���r��xw�4�3M�$�_"x)��E?yt�w��'��m���4��K��@�
y���(�r��PQ��O,�v��.�����!}�����b���
[��_�1�n_��~B��j�����ό��X��1x��w$f��LM��G��X��Ux��L,����j�a�^�o�JՓ��(G��!d�o�㙓.���p�6��4�|��3R����=	߁9����?��L�\�%�KJ���T��]�,�k���9��-~&o]����^x�%���b��x*v��ݺ��L#��hb�zQo�m�ª�"���[��oq�l�a�����;���e���p�.�7�ڃa~C(S���Vޠ�?Xxr���K=Y�eN�C�
��Lt7�����]���
�88��m�Jm>Ko�����d���U����-�)�Q ��<�p�S;-�~S��O�.,�c	��k&�� Ë������X�'rT��[[|c��n���'2�mK�!���qeL������SOg����S▌z�n9w��?�/���wYK��Hbh�&�׺+]�E�mж�#�u�.����d���zi�&�'�N2��� ĮC��}c�ۑh�0!�r�ڇ��O��T0�ӿ�Zٱ�Qzn8��/]Q�zE��2��oe	���>;���v�������\.ˬw<H��O��`�U7X�]�d����i��7����<n��'�l͛�#�j��E첩w�ȅ�U=@~q���x�t'8�ϻ��ÍB(� ��оm�x�Z}C����b��cGȷ�S��ޥ2�Kq�Z2�o��ze��_(�m����K=*�mI)W
�o:X�����n����)�~0�b޶�>����
'^�1}��ݓ4#�o�Q��v^�`��8�	�'�6�E��uӌ�p�B��Z�J�.��zFի�2�AN���\�H+�i!��n�Q���w�*�v?�;�h<E�u�jN)��MJ���q?Zu#�n��D/���Rҹ�4cQ`<cW�f%Gug[\G;�������4{B�p�Yű��r�����ߧ��܇hxP}l��/��t���^��)O{�uK�!(4M:u�zP�t/�w���`V��N���?��߆l'D_b�5�?��L��h�)mfe���q�������A�;0�
3P=����F8�8c�sT�2`A|�%�M���*��Q����H[J��z��6�h�^�|Ċ��lb%��D}1䙢���	�O?�&WM����">�w���N��k��0��	�xYP(��{qK�������?�M�_�H�w�!�g$v��.mv���&���lc�B8��&hm���E��6֨���Q�:�E�VNOZ��l�K C@W��)	agP�Σ>�l9��q��W�e�����I'<�iyM�>���r�J��cDڊ�� ���2�b�NZ�����*��u�����O���,�m7�J9�	���L�ˀ+����o".҅����A���)�u,�RY�\i��T"@�MI��iZ��j�7�d�,������Sn����+M���pV-�.1�G�i-�dГJ��J�Eˡ��yr]�by����E����~�>�*)$������T�ϐ�'������qcg�͖%w}������(2L��[i���e$��D�6]��O/a'�Ed�F�iC��S.�,pNJ>#fH������R��𶽟off`E��JH�<8Wv����'>@&��z�#
��w�v�K�(U�b�3uV�dΊ�0)(A$7�`�M�1Π�S�� *J��(�v~�.I�Q�i�#LN]�*Jh�N)�=�1��٦�u����L�	%)���y�W:�7	ٻ�Ͼ�6�G4��f�s�����9������%�-o�7?�1�.=<Ȅ�,��l:vQ&/ӟ �j9�v�q.��RSd�o��c��
�V����М�S��R����Mb��;k��P%j!��&���{��Da���܆�`�l�XZ@Q+ �s���߻�1���Lz�c��.3L��P�կ_	in�s�<}����Ȁ�~���as�����-�]���~Lv�
^��}�Nx�=�H�T#��X�^|�}9�C+��Ë��Q�
���	P�y�y����y��́)�R��Z�W*&��?�=Q�t��7���^���.4�E��Nnm"V�l~�Ͷ�Ew�O�B�O�F`�� ">T�8*Ƀ���5�pO0f�MBtn� ���q�N��q?�P��^�^P�,~�z�Xb�7B�﷝76z�6�|7Z�%Zb��-QJֱ]�w�^�Y�+̇y��̓��a����GX�BƝ]Ϡdt-��P�'s�������]A�	�w�����N+'�iWI��Ա�����H�U ͜�������썥[s*pٮ�C�2�����"���z)�[lͱo�
4W���s������eUE(e�ӤO�}�	H��Љ�W��iH�:OS�`֥�"m�_��|�N�:�E�ɏ�@��s9n�I`�B���5�|iS9H�4�q�C���<���|�RSϻ��3��V13�e�}��|(��?�(g>	�>��.i���6U{�ê��{-�Jyг'�>J ��Yb����]]6�:���,�*A��(s��J�N6y�.�!��A%�!v�?���8	�=��.3>�A ���+Iꀒ!�N8��{o���&� �y&�z�Ll{E���5C�րK��0��)�Ùހۙ���ҵ<�:���È�o������x�[����x�ؾf��0l�C;������"�,�M8KM��P�*��2�%�v�Ǿ+�R
Pm��⌥aJ�*@�3���eeG"�xAzx��n? ��1�^p��ʵ4U�f��k��޼��?nħevn��z�Pݲ�U)���K�N���g�;h2��N$���$��m�dKa����y�C!<L�]@?c�����k_� �_o��N^�ଔub�2iv���t�P�v��%`��.>҆7$�J`G��&�;��k�����h�z�����_���0���'�JC]I�<&a�[����P�̓i������fE��2Y"��e&{���:8"	����\&i�Qb�SV/�-�k�=ʉU~V�bp��}�(�B�����3�'"ƯK�g?��������4��nȈ)�ԯ�kUs�ڠ;�6�]�Ge��Zs��S΁Ψ
_7���#=�acb��X!�03ۄ�q��pꂁ�ܹw>o�գ����Y�أ-��%�Sra�G ��0���ؒ��3�����w/ɼ:�N�vjQ0xpO�=�����}z�[��f>�L��_�����VXh���0�9��ɨ�����v�q��_�[��Y	�k��	�9��#�"��3mU��k��B��-G�1�'&�[�W�iӭ�գ��j�挣6��/9�x���L���X��P�?�&$ԀnR!Apb-�����#QIgn<Y�T�2h�!2�o(��Y�PZ͙�"9��H�Ni1��a�|��jn��Gڌ�%����̣�4p W�z��W*���9;���Iu?�I�� ��A�r�?~2�t�7~�u�ǌ�`��������ʃ��X�����蜢��ɤ&/;f7�+�ymV��o��-$@�QO�.- ���_��=|y�oK�-yD&�uf/ZUN|�/�>����ԅ�,���C2�{�`��[��v۸�CC�M�_}��2�G/�ݿa�"�3���r>b#8�}I���mx���ʆ�#��_ƦD_!�:�UD@�sOGkE��C��&Iqb�ȷ`Bq2 ^`oC��r�S	c���Yd���\6<(wp$���➵�m8r�ћq��&�o9ҙf�L�a���r�a�[�劊gv�t��p�+w���uF��E���(�Rn������k���*\�>���}w1N�4m���@�m67>��y����{=����55]q�i$���H��-j�����D�oQ����D��Qj�n�f�p~�� {HN��'�!O_¹t۷�pr�����]�Í���"0�|�Ò.���x�wR���9�h]�����L�!L��Hv7"<N��)�P}L#�)�ǝ�� �5��,�O���z :#4_�[�������_�@9|,>pʌ	�09�H�v��e��#'�w����l�T��W-�^��:+�Ж��f��
h�[�M��e�A(d��P� ��������<� ��.��L4� K�+`MX�+����,�]���.fz�/���#�a��spFBZ��a��-R��6�Q��i\q�W4K;0M�*Gq
?� u��U5��ф��|���2̫c4��C����һ��ׂ���5
z�6eg곻%!ϭ��%Xd��;vc����C�ى��4��P�685f���f/�}M1`�Cg!@ȑ�=#���9i��f�>�'7m���)��mIԡ�&[ѕq3
S�$J�c,.���� `]�b���!r�3M��9�r^����ZW�~��R��e�-�S6�σ'�*Q�+l�#n��ڝ8��4I�RM��`Ā��u��&�����R��5���;aH����g���!r?�������p�D��	:.;���#���,aV4�
��a��h�fYb�֪�����Z����K�?-�Ύ��$�:�`U\���۲�ݩǲ;xGL�.M�� ��̅�������GZ��AK�:O��id�z�.�_�;xK����w����jXS88�M�������y��y3����5:}�3��8o5X燞TX�?�zX��+3�����6f���Fۜ��#�R	�(H�Ieb�I4R�di��5������0���p��t��`��o�'����8�t�|�t��L�З�|�`>�L!O�K^���=ð�����Hl���ƛ��N�IOs�#���k>�V�a�q��d���d�&r҇a��M�Wj����ꐛ��4�K¤&8��~��h�;UXU�	"-�\��؅�\�޻�K:To�4Ⲇ?b�q�j@�M(�%'��v���
d��0���η�/�ͽ���X,��k�؁�M�u��VP|����X�>�3�V�MG��;IaWD�<T�,-Go�΅���N)�����5��P����m���&�p.��h5�RI��㦋:�L�����Q\5d�u~ߤL�?([ ������n(@�S�J���Gz0P�h���g_얖�)��#�#�ߐm^"|:!)�zL˸�F�{��{3q��|G�&P������ &����ŷ�JGL���-�>ꗮa��}���{a)�N�EZ�-�i�q�	�J7O"m�/m
��.~���i֔A��c�~�wtf�;�Z=�����(lޣkjNqG��w/��S�F^��]��	?�Þ�ۉHC@p����5��~��۲���m;�+:4��dh��`�����r�o;W�@C�c�����׺�$k�0f��`*r��L���^<j�����)n G��>}&���<|g�'�3o��6�2�S�,�I~���<�c@�ɡг�;�i`i����c�_�x%Q:3mZN<G	�z_�l(n��;��Q������R!k���l�r��D�*���M��w��C`���nm*��T�\�J���`|��æ�r[�߃����œQ:!���b&�	�;�C�5�t$��A���W�6t�#HH2�E�����D��Z�۫Bm��U�[d=3D���!2�:��7��u�]<���� ���'�{� й��O�kc҂�mx	�̘�|U�6޸��d[�"Ѥ�.p�X
U�Yj��G��~K�I�Z�K+]�� |	��kݶp�z����^y۔�"=a�KA:J�NBq_��.iI-1q���''����ZJ�{���"�M��VKPTĞ��I�
4���w�����EĖ����<:�ּ�$��E�kp��t���"{g�!��Љ�8�-��{ֱ�_��@&P��e�ε_'!��?9#�>��W�n}�?�޶��-�T@(�����^���/7�ꊫ4��zY���(*jXV�ˍ���{
vٳӿ�Ν��[���+�ٷ��ϧtN�m��y�;ȓf&R@�E�	jj[j����8�L9fi��fEt�]i��Ͷ	 .��� 5���WmX�����3�G�]����54t�� �v�iH���\�͚ˁdx�?�I)L�<���FL�V�(�W�X����*��o��!��z��?6,�U���8/A�s�ͫ�.�aU�-�9�~�ᱴ��(�	W�������?�^�U_��J6t}�6�7���p
13;�HMx�1�HRE���Ǖ5��Tk�2)y2C���~q4�P�2��F#\m�Љz�#_«f`��QP���s��R��q+J_�ٞj�..W��q�M�C���C|�σYФi9�E�6������h��7½L�z^�[�I�њ��B@<��U̗�{E��).�����.p�|΅���l�V�̄ȱS�G93��*>�A�B���[�t�j_ ,��Z鉓��$����Cؐ��&��`X��C�7�B�h{?��^�?k�<3&�۱	8cN;|�o{�xp���q�~��-�D����{��s ���ͥ)­����c��_xV2���O�X���U�w���g-|亴��lNc˚��{?"_!�zѝ^wt��.��-�qS�g=F�8��0v�gr�e�7Ɉ%1�ZՙU���W����o|:�F��8�Rx$��Y�}��d-�V��;�z�
�T=�0ք���YZ8��;�����&0ܝ�i:O���r�\{�T�#�i�����!n�����2��A=����ཉ#�
D���N��5���@��As|���6�R��R�Y0�$mc��ɦ����A����"��	Չ��C�_B`�v7��'DVy��2���P0���͏��Q�S�+����-��50�3��'ɤ�|)mh�/B7E��o~����e���*L�Ӎ��[���5x=��<àu�L-� UEEkWv/�����2Es�מ�8��������]���tx�5�Rd^˽~?���KT�#8i=}zc�%sN�nLe��<2��HS�AM�K/�AKL7���~��7��J�������i~X)������z ��1>� ���� �9nv�x�`VX�7(R�PP���.)�7�!��+7'��6x��l ?i���Du��o�,�TW�F�ކ��� �<����5:��X�V`����!���lO�F"�%�����Q�2_0(���[���]�݈~�?�p�$���ȼ�R�A���1Z���M�Dp�Ӓ�#���ip��ot���BF�"��D ������.��N�����B����qI��+ ��&{��9�A�����zR����	�Ĉr� ��f���%�+^z, ,}ы�	,�&�7��!3�h̤^L�eT��������``3M�ʒ�����żEPh#6�Ja|K�>()�b��;8� �l���P\�,���;��[�v���+U���6�2 ������z?�b|^���<��ԗ��o֙�O�ar�л};�p4荗3�Km�
;x�?t�0��'r1o��m�f̓r}ok�7xu���7*I
@��pں�U�R.k�T#�
���u6���	��11և
��(�&���FS�����}Vr��-Ұ뺳p#~d�q�����̨����o}���.iWY�=5iH,�8��֩��g�Tr+L-]���ׂ��l�5ˮ/�%"��[:�.~U[\��v��K�Ru�KǘL�Le@�J�嶽�p4�����K3��n8aϣ��Hk�f<� �R���B��u�'bFgR�{
FoKP�	@�u$R��и�����H�G��c	�P\K�|�yv:\��3�L㯐 c�F0<��5��
�*�L�Ϗގep���{�{��`6�c8��)<��L�$K��_�����E�9�Y���X�`�&�	�~|�������qFM����C��ت ?*��e9˕+�^�7'L���]��N����g������+����Ix�|�I�:
�2�Ꮿ���o��V�:�l'm��ǭ48A�Z�r�نr��6=�(QN0�SMg媛g׵�\�����p��m�?4�A����X]RX]i��^�!J���&���HsK~k*��7t~��! �����ʇ$O��Q>5%���c~-t0�;Or�B�f
������"*�2��������bT�W�d��w���`Z��:�қe�S�ȐŶ�U���}�8Fh�$B9�E�tţ����G	^���yjK�_/42:�z/˥��c�����Һ���5q  �\@�������nx��T�fE�̷�r�&2��v����p�e��~��F�����n��J�O���e-��n�Sn8Z$,��Q3(��S;�?Pj�,�=��Fe*6��PI������Sve{���zޏ��%�A�@kHFBBU�e"(0|�F��&AoҢ��.;�<���s�Yz�/r�Ƴ�NQ���As+ɸii����PeOY�5�C��B0ɐ!G粰�D��u '#��2fҀ��GE�Ʉm���E����`�`w�{�_�wO�6����gt��nI���?+D�7��`�5gw�v�5P=z��3��o��pTD��3K��y�;ْ]��I�����T��r[#�ڍۚ���pg���b�'r�߲&��M=g_�2�R�Vq-B�Ӱ�z�`IB��-�~��J�C����}�>�f��x���AZn���h;�`�}������1V�g�.#��|"%M����E�ݿ���b�l�Hlا_���D��5Ӿu�Yų�4;Q&��!�� 4�{Kgoe'Ƴw�t8?|�R�����}�ߡ�kU	}x�[K��- z�z��d��6�G�PE8�λ7j���V��sq�>bkK:�Ԟ�59�M$���j��K��`ؿ����i1���@��yvn�^���K��P�w��� Ұ�s��;}�1=<
�p�� ����s��mQ�,�?�?�L�e���2���l���#�זݫ������6K�l�R���!t�]7�X����ʧ-{Y`�5��7�.�{,���f�zy:���EEY��زn9+
����)s�~�E�F�O��hlqw�#Q����Ʈ����j���!>O;�"/f�(1	�7$�s���wf
S�x�<Ch�b%���"�6M�Og
w��ui=(��P���ݜ�!��}��x��r���ʓ����w�<�h��)^jadTi��3��~�lf?Xp�C��H,���H�oȩ61!���$X�1'f�'G1����F��9~�l-wDNj���B����:3����m����)k9��O�ɕq���ꃯ���ʓ��6�k�ڷݩ;�8ZB\?&�>���˔H�w���P�c	QO�ᵙ%�5��!XD歯����\,�֝�]i�RQ�1}r��t\��]����(rf�X�O����D6�@93\�Y� ��:�[~�T2/�m�nIL3Ȃ�a5gS�뭹�����VT�p�?W��˥2��X�1�SC�ਊ�����kD�z��Yw���D:�+k�����fh�Nn�zPϕ��H�	Z�uEщ�`�	�F�����6�y�ط����&�=RW�VZ��C���ę�_�-)!6�4��Vz������M�i5�����znsi��8���N�� �����bbw�,�*��~�ͅ	6��	u�[abL�Z�&C�����o��UZ��R�S&��e��x�����KC+H�Is=��7�{�`L-ǿ�6	i�����L�R�C�x޽'�us� l��M����'nK���x����g�W��7"�[g�\(���f=��K��ӧ�H�IK��#�%���t�Wt�ܛ��S�����3��>��BC�E2� /��t��nw��X�Z/ۣ��}�5��>~Q�s�=nX����g��6�&����u3xH��l�2T.$��46$ړ1�����*����wL<���������u+�F=�r�0~=0�&AHr:)�	��Ff�o0�wKZ�}��K$hJ�Q�QK����r�Uu�E��F:e����?7�-��j[�����f��o��:��]~[ζ)j<�~']p-Z�(�֘Ei��ս��;Or�sb�]������������f�bW����Ԃ�R�u+��C�7��k;��+�|�$�E�`7�}%��x�]�_"�R����i�T�f�P�������6��eG�H4<ĸ�n����m�^����K �fdxld+V��|.�#B���>6��Hu�];��PJ�"���.�<j�#/u���M��&�u+���jٷ�[�ѷ�)US1ʼ��c�i	37��E��B�,��."��EZ4�F(�u�~�]���=
��Cq���-t�<�<�vD�+j)�q���o_�Y|�i�Ueu��w�]�|JT����(��1��w����I���_.��/��b�+�RϳRu1��p�H�v����$b�IP� ���Hhn�,)����燘`�������	Y+aB�GT@a����N#�Q[W����vST��@P� X}ٞ2���0M ��8����L(���iԸ8?{���Jt�,����F�n\N���zX(a'[S���mɛ�m��w�����D��������>�O��<	V$�nqQ�b��Z7O�;1#�H��7z�*Z�dچk򳊭�Y����~��A
���c>в��E��j�'u��w����@Z���(U�e&R"u�ߏca�Z!����P������DTnۜ罅\����M�@��O�@�]D������@���7����x������	6���^��YN�����
De��k��! �8۫J�8�AZġ	���r/��_�l�U��wGjV��@��*{��΅(���C��T8W(�U��Va&�28�a����R2,y�dD�R�R5�^G��/�{�����\by.It����̿��m�_vc;�F��N���y	��iX_}7�k4��vj��|���q��n硤��C�o��]�i�#B�{e�uܐ��F-��>���X���4����.p�W��z����ҪN\���PI�H㈍:�r5��xzg�4T��Iy���VŞ.Mz��3�݊�\��d��A���R��m��=��]S��{�ת�}�!&�fr��_� Ts����Egd���9�B���os��8�%@�D����#h,1�K()ҹ��W�����I�u�*%�u����V�<v/  *�i��>T;nj͡.J�'B��-i1�����' .�yuB��(��b?���Uq�"L���{v��{�MHͺ�������Oȇ`E�P� h��ݮZ����w{��1w�O�6q6���`j�6�D�˻A�9����0��m݈�J4�-��幦��4&/�ѫh
�6�?n��'c�'�(�=��ZZ"̍?o���~mk�a�ǫ�~����K;G:�w����!o��f��2��Z�7FΘ��m����q��J'�D�ϥ�z��|�[tѱ�x�%�{��Iy\��Q�a8��Oˠ�aM;���n��>�|������8��f�%��fjd��ȍ6�@	����\����kw=+�d���W�9R%��q���]>��)����
B�e�e�ou6���`�6�\Yٵ-)�Ew&�ס7QP�r��Ch���a{"�?og��ɯ�>�`��/���_�^|��:P�8�8��(~N����;�I7;�w�ɖ����*/���]��t,���|n�,�p?F9�Sx"���K5�0Q�6�$�B�Y�T>�nˣ�U�d�Z>v��0@,�b���k�Sr?�AƏn�=��y��gwFy���#e��{zW�EAap��w&�I ×�=g���s��곆	(��H�ҊT]ؾE��I�3�#|�q"O���JM��U�5��@��'�6��I�=�?�����.H3����T]y<f F��g,�'y�))�����9���c ^&��5�Z���g���&�x=I��M��K2��4W��yq	OㄨO��
�9����qP���ʴЕ�r|�^J����`i���Mp#��}�%����{�$#o�8\ fF6Go���~��bba����!����5zT(�3,ٺ��/u�;�DYR���#Fl�*��e��Z�rя]�R��0ަ��ݼ�Fk��*��o
�K0��0yM���Qp%�#�`J�M�ן��l��@t��HL�(o�z-�1+~���Ԕ���g��7�ڦ薓���CU��j��T�gL�C�� �/���0t-l����xy�ϣO��D���$.����>f��d�[�^x ��O�P�F;-�HNI2�����������ע�L��i\�'r{h�OJ�d�A@��cE׺�
/J�aM��%����w��Q-�w�����tyF�T�8��Ք�UI W��f��poa�S�T�E2�㺀6�h�/q�s�~���9�0���f��IU�������U��gh^CIo�۵b���u0�Б�
��y��^���#�3�=7kt�u�����}0GL�Y�ɦ�?5�����)��~'�|=]�}>�@Y�h���\!�Ji���S;G�+�k�X2���?�Y�	\Z`o#�֝h��\�;�2ώ���Q}����':5��K��R����U-@��=�^�t����J�:�<`c�I}��g�����)V��8���������T����2u%_e�R0ÑpWͧ  b`�t��ö3�U�����@$f>i�wGƾ�L�q�7.�]Mi�<�����hQK� |�:���5<K��:qEW��Կ�$,;��rq�@��w�O��Ok4�k��z�u��:���
����U�a��E%���8�,^)'L����K���:7�V/�q@Qxf�ٝ���[j2F�Yu�'M>k��%N��գ'ߵM�ԃ37?i?�F��zg����]aY�[E�U*�{�=+D`ь���fV^>��X����'n��zee��Vٌy}�
�����+��0j6U�b�a��C0u�#�U�����n���.�+�kDV&~3�(_�����q~n�6�3E���Cg��i��c�`�l��+�3ٜ�8G�a�$�8��ċV.[���$[�cOڈ�j��X
_Z!��F5߻���u���B��cQp�O_e��qE�] 5�-��]+z'��-|�j�&1�A�9L�1(��Z��E��{��A���Q��ޙqа�	�M9����V��KHv����V�o��ۡ��=�����4�V#G��c�Ơ~v^̓���K��Ŧ�	�(�����	v8L����!`�cJ��pMs#X!WlB��W�p0H��������;�e=����)���X3hy��u�&^���I��Fa��~���r�8\񃏯F�;�b��ᗒ�c���SgGڧ@�sDh�D�e�kQ\G�j��pG+�i�b�(�^�L�)m�F���@s1����h�"���B+85�/�g�ԥ3���A�u�ԶW���֐�FZצ�6E9U.-%��ߊ�>a�ŃF�X��տ5ض����v�+�/_p��~�+���w6�~�M�	m�|���C��ݴ�7�������ޟKǞ!�����L��.���m1A9)��R�9.e^3':�]�	�;-J��+�^��{N�����h�H/��6&8:8�8�Q@5՗3��VH�g@�L6�Q^�F��ѩ�YyDi���	D�ow<S�7I���l��r"� �J|V��y���h�vI"�����:f�@;�('*\*���dNOܳ_[dY��ӝaAm�cVk6��+c��e��� �i���X`�x��] �&��db�P�����ڳq'ƌ�Z��R,��9kw.�;�q̚]�()��c��<��A�	�`�TB��-࠳�e�Z,�Ӛx��4�$ڥ����cw�/P���d]�lZB����O����u�lY:�("�$��
]�^B��|��X`s�YM�s��DJD(º�I���^���1R�������<���nc	:��IaA��Im5ݥ�"7��m��̡��f"��<xN���@���8p�
0I�������ev�ǔ�7m��������%�
����Tl�u����q�[�Z�`�u��[��(̐�_$�OjL��y����B����:�յ����`��f��	n�A9v�b� ���ď��RU H�
�1)зڸ}�4rC%r�mZSOr�77���p�2�{��:LQ�cŊj&;��PL�3�χd@LZY|XJ'�)�J��"6Ʒ�c:K}�_���8,d�U�U��VJ��n �GƊ$d�:��8�G'h1��L�D�!G�Y�	�	ߞ�¢� ���=2����/d7��,��
����0'�W�.�[�X����0]wIo���h��!h&���1�[�2�.Ҵ;��]�I69eE9Om��0���{�M6��P�0�1�#D��>S��`G��c����T��Hz�x}��A�oxy��~�L��.43��Z$Vb:8K������FJ�m�g��#����ο�'�@�<��HA��p��<,�a2�H���d�)�t�����=�?R�_J�N�H�3�x �E'�7��u��7>e�z-ڜ�}������X,6K!���V%t�v�Ƃ�Ñ�j~U����-������}~�����j�s[	� `��y��TTk'�C�?���1F����,�-Q_�)	�_gJ(��)��Z�V�X��oC��D�
wK�_Hs\	�̾��w���-.0o
�l�n���Z'|�Z]Y@X&��T��M 2�����*�B�ͽ�[M�Z�R0��&��-�)�P��8�*ٰ	x������?�����a�'7��,��W���{����]f��f��m��dy��|ևPm��x{܂tiĦ�)f�,�l&�U-O��c �P�K�x�F�@~��F�r3�����|�prC�۳!-�T���D�߻k�ْ�M̈�F1��MD	��r\�"�rlB�âwNg~�Oڕ78�uu��Sۢ�?�$?0 -��/��"u�1y"O#e#��)(���-�~8zx>��c��K������O,7��o�#F�Qn~x/Y����<|�w��\C͚�#A�E�V�ZnA3Q���|Ud��x#����V�}�|Mϐ%@��B�V���O8��W`�\O�A�$���+��e�",�� �d�����1Uʾ���km'0����Κ���ECv ���tBO�)�M*�M�
�M
�����# ���[A�ӝ������'j,��Fް���2x���W�w��2������Ԕ!��v=��5��W�U,��,l����KM��"!�OL�Sd*(:1`Z�N'���dܵJN��S�}�/�ܺ(+�&T(UHN�©h�r�vck�}�SL-��6(�O�X�4�Guw[e�Z~�2R��A�/+W�x�P��9VN��L�~�Eb����c�˱+	֟�_��	�v��,��[���NyBrЭi.jȓ�)���@(?�5.w��U�6����wZ~#�O����T(��}����������}_�#m��=�?���1BǸ�1k��U����F� 侂O���n��&�
5��� �4��١g���gm�#f<�.!t�2{ ,rhI,-���V��=k��yk�O ������H*n�]�J]�Q}���n������I���6��ի;0'��������Wn�ͅ$�<��TmS�I��\������:c,�E�od�<a��*"�j���93&"�� �d���x��P@&��N9���k#@έ6{������W3�`B��빚�xխp�ze
R�h�Z���\kB���Rj��;VL���ό�M���52l�w�٫x����I�>ИY5S��|���J�>��l<��ֱ�|˿��{n��Ur{�aL��MK�ٛz�l�@��eDI\Mp�Y�&{�	J7��Y���Mz0U���oi��><4�;�!�����/�VM�*�{�Ij�㓚Z���'x"W}o��.:T�����-4��g��|�aE�vmhpB�&�i�xu	�f�f4)�%�	]���������Y�{��jZj�^����t�J�sx� |�b��V�"���B�\>�z%�Y/����y5Ec(�%�p�M(^��u|G����B$ɜMn�*}��-�t�26�(2�e�fmb�
F�ftbF�ZF�pB������%���K��y�S�`!���W�p��2�gF�	+&�+��Í�k�l��@��uT0 G������#7�מ�pq�N.��=T�ZtA��K`B�W󂜄(4��E+��Y0�I�"-�.���Nw��z��6{W���hnM"�^O	*}�6���!)ؿ��m��(F& ��q�b�M��J�6��:�
�����J⿞�������hS��_i�m)BL�]]�-�ִ/����A&����~�j}�h����LI�\�3(���p�=�r�#/��uR�?�C1z��yp�����W�Cu;��/t�l�ri���x��<4���K1p� _"3� =I����#��'�U�J��iF��c�9NJ�:E�[��.��Lۭ�����]���تA!~d�*.��� �$��~:gNx��8J����hf%_7aH�"ݐ1�\8�ӷϧ*2��[T���VP��{�̊W6	>�,=�п�Y�i@��f���֙Z#�2��B,����O��-�px��M?�g���m8�����|���m�߉�Ǻ��?�9�U\iU��hӲy�FaI�)۾�n���Rx��,|��,6���f��g�? �	��Tvx�����c�Ͳ]#W*�yi�o?`�EK�+�u��A�Pr�Y \.���<�����!,Z�=R{���D՜x��y>�Pj�m\�	�]��.�#�b���ޠ����;�^ʡ���*�'��$;o�@HE�v"�ձx�N	�n��>�ڮ�V;�:��GA.M5���ӷ�+����z^S�+.��xX�'�^�����2#2�Wjm���e�bS3�&�}Z(��F z$o7h�����Eq���c��6��L�@�h졙�(�!�����][5��<�4����	��i�v*Ҫi�eUT'�Y��ST�!�#Ov���a6VRa��hE�!��ͅM���Ӊ�J)��CH�U�Xe��W�� �e�S���v�:DcQ�����m��xzw�D�6�O!?��|(��&\=SY+Y��M����]����u�=7]�M>�+��z��f��	�H^����;h�m	g<y#��8��mW�[*����R8P����0��i���N�bi���é��O��Z5��Rl3 �=ؼ�Gǐ��'�d��3:�I������=5"��&�M��o���j0o�6�˴O;�����>��,��~o�.�|2��8����ʭHu T��4#^�n6��N����r�>�:�M�<�J�f8	�a��������f�e|��;�������@��-�Xݴ�8�˩0�����Y��m��t}���P^>��E���<3�@;`[ �M?���F� �G��]�Sd2Dϊ1��W4�>2�h.��+�vOaQPQ�
�;��Q��R1YzP�Y�|����ܞ'Bɧ�?�)}yVP3<�e�p� iV|�dń�������$H�Iu4o�{�ƫ���u�tx��q���H�nWv�=Y���ІX�fƶ>vƻm܉��B���_!���D7�]o|=��V�TQ]t�V���#��������L�V	�\���l6�f�XH9Ʃ<����q�X�0�,��H
V�xb�`xn/J�^�}�f�I�)n�FZe�ېh����a]c�
np-��͛�	�RIPfKױ��/���!��{r|�{��wK�wo��i<��#Y�6��Y��Y�U�\ֱ.Ｕ)��Z&IS���Np�F����%a�|q��^��u"@��ŢA�t!Hߌ��P��5��n��G��L�@�����K����0a��@�"��7ݖ-���	qo���Ł�[1�!�9D]�^�6���_�ޘg�`�o^��u����C���>X�E�%�o�#�]�f�H�G2��B\�r�>� !ܖI��M��Ȋĉˎ#���Gfcc�F�t�f�?$CR�eXГӣ�4s��[�;S���ˮUR=���y�kĪ�$� �:V:�K��?�>�L�d�1Av��~'��6�}�����M-S�>P
!�!j
�o*p������w��1�	�?EȾW������Ng����Y)��!�_g@���J�6� �)��)�Oq�����O��\ʭ�N�r;J2L�����E�r�q��-c8���C��Y7��X�Y�H�}?���w���ȍ�.b���M>� �d�L�S��?��N<�p��Q�94�� 1崥=���J�i/�i8�@� ��8_p���ũ������y�51��;Y�P�w3�9 >~EZL�P�"I���)T�9��uAl�>q�^M#K���ܱ�f �����k��!j���p����%�b[�Sa잸R��ʦ�f��z���A�'�X���IE*�O���e�K�|�ݬ��n�#�-���Qچ��k[��[>W?LW7m�?ɘԎ����ִ��k��V:U�w�ৢ�k @hq�9s6��mzM����,U�.@��1kv⚬���2{9��o��{S(.}��hd��?��o i_~��V����^ԩG;�P��V^=�\T�S٧�ja��q&	H�?���ޟ��+�"�t��y?�����D���'t�,0X���������9?��rjӜ��`�F�%\���_	�6�V�������;�ϘC����Z7��?�P7�慵���Kŝ�Wi��p���m���^vO�p�ꯋ�̒�s�eFD*���"�h�l[�]ωQ l5d&�	�a!f�l�:t�j�3_������Y�
R-�%0D����
�B���,TPԓ��R�,cQs��:�sX���Oq��g]��o܌>*(sHi�shﾹ�m�uФ$T��%�'��%�k���̡Y���8�ٿ��q�������Qd��&`1C!�e�<ɘQ�����F7�(��Dq{y���qB]\�8%�.�1;maW�F�S2�k#iG^w�\�gY�o9��eb�=#�j~֛�0�.�x8�	�^�ޒ�wq'q��(&�0�N� �
I�t�y�G�Lc4��/�)��q��w��ka�z���^��ب�zEe�@��W��X9����y~-;�ג��^�f������<Ϭ��|�|;�����Ji� �+�ḣ����5��#`m`������1�7k���F6y��x?���f�/zA�s�@�U�ކy-Mad�dnf��qz�����t�ȿ눔�����jje�9wǃ)4��Kll�0XkF����D�&V�m[{뇃�-x7��8�,s�/������$��y�AM����e.��l,i���1Q|�0l��i33���τ������5����i� ���G�7|9��px@l�%"C�(��s "b��˵C��g�o�aS�3����`�hMb��lq��O(>,!�ş���������sg���(��r�����7�c�ɤ�}^n�&��н����C�,Ay0�sSԵ��V������V�n"	'�O؍�J)�$֫#fp	v�h�[r�#�
�?}��ҋ���7���L�>�?�s]8d?f2w-�QP�泯�,�A��`����F
Z*���b�PK�.<n�����|���?�Nj��}�*h}Ԕ�Z�g�l��X�}�4�l����r���^�LUd up�q�E�[�D(�ћ��|�]��yP,��߃��(���q�g�S�2���Lw�������iX<?�`q����~ σ�*Tu.Z�99u���l���E���#��48d�M+���E���*qC����g
��V3i���I�G�U���q�`��Ձ�����%!�&���lz\�����H9��-�J)�B��"}��9`���9ZBm^��4hh}Hrz_���-#U��Oc��6�oOŧe�wC�g�Xג1;�p��ߣ���7��<��=/aX��=H%��5�[��	vmF]>'���~��+��j�~�yJ_j�ʁ��@<7�w0�
T�~��^X���M�TV��G8�8���e}gs�[7uKdɽ�������b���ef}�'��XD'3��B�<Y#�8U1�(�p���>���ߡە�Ev�j��?�P�W�r|l�oĥfq�]
u�|�|�n�нyOF�6ry�#��H�*ʧP����pTT�W�~p���S���u�1g@p��T���<�̻�����b0��g�8�Bb����6�5���Jk�~�[��t~�9�=���5��|Rh�^���"X�Y���l��A8��Ǭ�;���5w��j��e~����	�^��E�>����wU��[Ǒh�6)��֛�a~���:��./��L]a���p-@G"&V��=Mƭe<�r�Ĕe.�1��Ŋ�KUM�-������-O`P�[%|@�e2�`��q.D_���J ��+����`��b�$��������bЯ�ỉw��ֿ+���F�B�|�g��F���l�Y��[�h|��Ubw����i4���ar��Y���z{��(�ˊfs���	��B�NX�{���� j�Rq�ٿ�����~��h�����`�3 Ltt���~�)x2tp�矜ȧ�UN����B�.��Ԙc�D)�s�I��P!KI�!G��bbq"��p�a쪒3��i�����%���u��V�<
���&���qޅ���X�Y����E��u��q�
�">�H4P�v>�=�ow�ji\9.l�6�����D�>,�5y��RL<i`�i֙+<c���_ �N ��zZ]n=�}�E{��[�ˇ!MjW�����cQ�!�{�R��L��;���=t��Ǖ\�Q��`��H�s=X�;�������'�C��O,=[�Ip ��]0c&(2���X��8�,�6���L�h����$���/M�'���a���W�ƅ���2��%��s���}rm���P�� ���W��*�f��Ys1����F�iΑ�~u|�Fc��2�8vw@Jj�ݗ:�H��K<}S5��˲��G�5����K�~����y����ѣ�"����d�y�L �iD]�җ`N�G��G٫����P�y#alt-%!7�PH��dFw�f+��p�����������i��+N�mh&�A7�O�*9Il��;�_��}�.��'OW=ʘ��E�>wА�1�c(����g��4;�ʌ��&���5y����
@����|ד�c���p��fכ
����l��0V��#�?R�m�i��M�,�C� 좷$� LQoe@&���32���9��X�<�w��2kr2��&���$�.'�`Lo��ߤŜ�=�N#��i�L��Qm����{��МťL����h9��b������]&�=9ё/����i&k5؛ߊ���h��59�G��Ĕa����"��∌r� ��q7p�4�Emr:��^�4м���u�V\�H��@H~?r�_����r�8r1W��[�/c����\��G�������M����Ŋ�����F���M����,0D��o�;e-�����B��c^y,N��b*M�E�u�ǎ8�K=�#��.T��s�:���+
w"��B�ƹ?<��T�U;RƲQ��c]^C��Z5M��XG����yj8y�XY�:/��e��I.�؊7�h1(���fԲn�eH~)|l@l�0��憍��~�"�V�F�y�,}��%�
/��3^5�$8�N;^�E� {��Z#_�J��9.5��霶e٢�f��S�Q����H�����E4s�G�Q�8�p�n�,���6Tv �L���G�!��K�K������nd^O�On�͑6Z�g;���'\sjJ���ƫ����B���,n<��D�#{���;�p�������ۀ��4�T�ۚs#�p�-v
�C��h>|��r��0ղ�8jb���(�K�h��R���a�MI_!k��S� �:n�
s�uIM���Z�dX7�e?�?z�39��`�UK�����P7���l�o�T���7��-#�2.e-BE����OF�H}.}��22�qxlj�h�%�M�--�%'jd�V����ֺ.��LՖ�)�ޫ��^�P����KCV��E��'�ɻڱF��eꮁ۶R��[�.�9����I����e0ф��h����[�02+�.�P��7hY��I�(���-�*�����̅�6�7:�J�Z>�a�3f�R�?u��J��9:&��`+�s*TC�6�*�NL� �X놙"yi�Eo�4��Y�y{�F�z��sA�rFd�CgV ŀ��i_憳ө������Л��? �c�O��GOeX.�a?�t��!���Y?e�l�~��MDA�v���*�W,�q�,�j_�g�+�WA�m��f�鰯N�,nX���6x��]��:u�0�t��v�.'���*Ą�[k=r��P6<o��`����/�5|��KDKE�_dS?��y�F� ä��嵶S��]��2���-!z�t��tl|��ӂ*�t{m=D������'E�X�Wd$��D}�j˲�NDФ��һ=�ۂ��1��7'_bs}���������2�A(�^m�4&Ȝ=�_�1;*��b�rx�.�������x��A�}���*/���Yl˓����L��-쉌�4a ���A��%}<H�.��:V�(�������`m��f�%�_naO���sG�k��S�+�w#z����νm?'p-��z&=�%t^6�&�z�4�`������WB!��nѭ����cI�?!D���G�)�F�)V��G�%�eryZ��*�i68���H��Z���%�|v	:�ɶ�#��Ͷ�xX��ƺ�AC��PȨ�t�y���L��L���yK�|%�6d�"^4[f�U4yd����H��,\	���*�fp+f��D��EZ�l���4bvy令2[=�J+���3ё�7�0c)<�`��rCI�C��$G��DR�k6}��6�������/�A�<����&����K]aJ���S��Bg�i:����m�{��:����m:@gg߳�Q��$q��v�L��M�ؕsorK��w�_�2�KRV�&rQ�"G_0��aK �E���{a;�I�.	[��*k�-�95f<'��.뫛Tr�����y�+�l'��,����q�{$9�0��Jy-�orz3��U38��{&���g��=����vn���w��@� ��S�A��*(�%��[SOZ�3$��T"�
jG����f�r5�Cj;�Q��{1��.�R�3cO
��}���^�Rv|���%���7b�%sl7gr�c��Kg�<澎�@�B���c�%�N�{�E��ϩ�Ɏ�9��J��:�Z�9�\C3��1K�i�Y��Ř�jK3���v�rL��\i��l[��'�u�~h�`�Y%�Y[�'����o����.۰x�>���Cl�����Ay9�ͪ�+�0��H0��a��ް[G����s����!8�CҾ�Yk�B�U�.5@� ��uϼ�^���>����L�������?��h��3E+QtPh�����$0�3�o���'0/�o�nO�w,�1���9&�Mn,4�xvԝW�q�S�K���9�g������re؀"��r��}{���Eܴ]{g�2Y;+َ�)�,7K�1%5�0BR�m���u!0����Y3$�k⌅�^H��J��J�ʑ��'�l�������z\���L��9���{���,�yy��ǜ�s�c�X���/�4�)�/,<�+��4|����n��W�P����^e��B�Z�y٪�m�r�o�I�"U������]5�Vr2g��ԟ��PF�^���._�3ޔ\��N�����ZLP�5�N���C#Bd��Y�n� �_۰jIA7�)�9��{�zna0��O
7����q��ʂV�=�eЯS�c.���;(�����;?�蒸8��<���U�E%I$Vr���eg�|ڲ��0V���d��W� 8��Rj,�#N�k�L��Dv�x�.�s7�V̭d�B���7zn*�e� W���{7��x���dz=q:U_q$-�/vu-�V_�M6p4m�<�@��R�������G��T+W�k	lE ��*������{����ϗ��h�@���.�h�̘��ڟ�)޹g�;=��ޕ���$E1O�#��s*�(�+uC��5H�
�b�b�q���$���t�4��\IO��|�T�
�_mh<��l��Z�s�o&�`����4bNrZM��F��� ��0�9O��Q�[���f''�c�����'C��2����\����ǀDO�FN�y��R�����8ª$vJ1����Q4G>�HdB,�e��o^�x2�<C������w5��ǈ�8�����?�*��JyB�k\���\Q��?q� �O�pNӪ��L���-��A�uY�'�{A�����R䌢b�q�*8'f}
����������D� zmC`Q7��4~��\<�Q+�
eI$0V�OE�nvG-��cW{���O+��QE�S����,I<'率�I��*\)��6V�;�El��9z�d%Q
R6�?�F�C������~�?n��l��*!#65*/�X�;�ƨ�,x�O
Faeq�N�k*��Z���-�0dO�*���j��ȍ�sd7��%����� I�0Ķ�G�����d�����){.�?��>�����"�Rh���~0#k�PP�o��.ם�9��&��.�#.�zٯ���J\)� >v��OϪD�����L@�H;EUq\u�vL�V�c�ղ:�T�gb��C?!�ᓵ^UJI�U��	����X���Bf����	W�R�Mp�a(���%��,ێզ�O�G�B�-b(��<{=�.��.�oX�n�VP9��}��Y�I櫝o6� d�u���-�~]*��K�l(b�) �(�мy*���eJ�~�V,2���3��%���}���������>�^*��Z(�\&~�n#�"�Y#���})�����~Qp��+3��i�'Z�V�!E��2j\YM
�s�q��8�R����%6E&-���I�#��U�͍.��L�a����i��q���K����`�P"T��)׆���ehd���\��-����Ȓ�]@ �1ԙ�>��J�;�`���a��?g�ыԣL��7Ut��HmH�;����NV�����&��Ԗ,+|� ���/���YXh����FI[�yW#��94��Wʃ0��!�7�1è��!MA�E�k��e��x�Ȍj�A��!�;�%�,OV44z[Aj���g�Q�9����ClhMH���R"��k�.h����ݔ��z���y�
�g�F'B���g"�r˂��~�/*H��T���rK��?^��P�/��u�{���r-��u*GJ�2��,`.f�58R�g��\
9s$J<��o���F� ����p��U��PFSZ��o0���[��[LMI���R�FJ�~���@�ģ�z�L,�����z'����0N���x�?"��a���������*�x��͸R]���B�5���אrbM/Q-�{R�-�:S`\��������r��<ʾpv���=�)&�n�U���f�>�Lv���+P{�M򈩻�؂�Kfd��\�A������l9o<�ݼ�f=Y�eZn��d����67&?[5��M��5}U��&#Jizԭ��j鈳�	��m�bL�T�B��vB�6嵈�0�#��^}ǔ" �-9f�z�4�V��E�3x)���J�aZ7�*8�V2�"s�_�5�+No�i�w�=%��	�
�.�7L3Q q<7��硡�����\sR�;�O7_V�hh��p��ק��Dh���!@g*��Me�|#/�A��di���n�T�_�ǋH�eB������Ҿ�.P۩�6�y����:�(���Z�V,"	h�@ƽY/F68�O�~w|�	M�0����(Ԅu���M�<�T�d�6N}	���	�5ƥ����.B�h��T`����?j��A�����ذr�փ����\6� ͧ��h���!A��}�	�K�y�0ݻ�RF����TV�r����*rS�XE�"��c�㝣�!��"�y��0Z7�[`j)���jġ8/�%��%Z�y��}KI�nߗS��؝,���m/���������m�3��e�_�MB	�`޸.���gl�{��zAR��x�x�����K�.*����zF�+��ajU�6���ϖ��?��/|W�X+u����E�V҉Jgb{����*�:����.S��U�}[��.�=��
�LR���`���;�u*Y	�Pf�`���D�%�<�77��lj��gDB�v�2|l�05�k�W7cV�}��J���N�x;�k�h"�Zݿ��x�A��~��4�Ix�@ɇ@�$W�0�|HI�߀u��H���c(�
���@�r D��=ִy�E>��]ƪ��w;āV�Y�ڦR�V
z���bu��M��~{C��g0��}iU�������&���{��I�8��-?��c�I����:�%l��:;&Y	;"efj��y?�"���l������p�"��Z�n����[M���*G�*���~��`��#���8��������P$����d,�n8�����M�*$��12�=C�L6hJe����ޚ��7^Hس��ƿt9�?�u���1
�Q�o%V�zo��&�n�	�@66(�ƺ������%�j(�Ь$Xŷڨ	ȎU�#62��q�p�c�YQl7�5i�ٖ[� ��w���=q
���p'��9PF�g�w���;�"�V�i��T47��������( 4�A_����H�
 ןD`��|:����[���nȧ���ih<�w&�� �iKk��;����:�؃�C�4`��g+���54L�>�^]M1�8��v �\�	<J�?,{���K0�Q�:�z���uP�imɟ�z��v&����i�f4�C\�k�ޛ�lrڨ
�?��Ah��.��7z���	(� �@R�f|��/�����ȭ�ğ��h�%�ٕ�5C��N�Z{Ã�m���,v=�)�vF�R� �3��{��kh�AIP�
�=�J��S�=5����v@e�"29Y��L	P�o`�����,.��������@+.
���.�ąm���v���Y.N��6NL�Z^O�1�Y#��uh����9�Ǜ!>�bR��*��7V0�{#h���f�Lx���-rE�����6���SB}U���J���O��._4�)D�
��?5%(��T������gV�%��+T�L�aw���ת����=}3,��7�xw2)9�|��>4K�R}�(��9U��B[D�\�������r�an�$����.�����:!�ZKB����JV��*DqO=�O+6�+li����s�D:��l������;W��')�fN�����!6�'y�����J��f�^�6-����vl�s�g�ɥ��}K N�����bb^��zt���������8 �E:����e�}�+�nw~Ƽt���V!4fSqc��3=��M�SH4�'�� "�W����Bp1b�r����4ӎ�쳣MĂ̠֟����Z��a8e"�<)T2�0�0'{q����2&��уWv��U���5ȶb�|�w�к,\݈�Q�="���^�[��d�၆!V�ۤ�'m��3$���^��ΫE�M7��܆�e�2*�W��Z>���:��]Ѓ{�U�v�`���&Y�����:	IL�*�0��TmD��c%xi��x���D���|mݢZ\��7�g�P$����tǂ�Sq}�O�:�T��|`�Z���c���-n�Pzo�9�[xq/���ޣ����J������\��T^�4B��RG�W,��D��`(>ԉ��q��'���Ƌ�� �+�I�,���<����� �bg��6����0�q{�x�o\�o��ſ�t]�]��32����J��`��4y��Si#7\0���1U&|!	X3�c/��J�+&��YM�g�r9��'�NS�����|��?��.9����r6(��Φ<��[�d�'�37�~�W=�>H����~>���_-爉�"������Һ��H�ݒ�m��4ϱ��I@�g#���FO-��$�f����͂W��/hU��=�d�5�{�c��bNpB���� �����Uz�6a��L��m��:�L��;i�q@���?!���U�3��"�0 ����&� k�_������K8��u���_B�c�@4l�1�� -�`��Nc�w��B�쀭�S��Guo&��d��I��c��&bq���#<�ŹUQ	`&��E+ѱy��*q�FNb�bM��B�į���`N��_3��C�駹Nm�yu�����C9��2j�[5h5(�/A
�;����ߺ>x�o�������l_[���O�O�"��9^�!�Mn�W�F���!��/ƚhUnq�j���pH\Fs�ўm+5��IA�9Xwq(-���lD�����q6�_y�p�f~��.^��0Q;@�I����e�}�|���C�:ŒV���(�'���5�y�V#����:�rw���f	z�ѩ����$h=�tɝ3ڛGȠF�� �: YU�a6gΈ}�Y�*�s�C���y�mViP��Ҏ`�*
ъ���z<(������_{#^,#%=�3~S�vCewJ֒��A/��z�'�d`���	ʅ8��҈��ֈ!7z&��!�횄��l"����ס7�������C,�d��7\v�E�*wkБv
��3�qY~�}�s���9���K�����W�v�n)��g:�����j6��&���$��f��`�@���D��	i%�@_���-w����߼h�٭��ɶ�0J�Hs��\T�C-��N�������E�%YLi��nN6h�.�_����Kr����E
��ad'���/t2�fH��mH���ҁ�Q�b����H���[����a��i�~ck�`q�b`E�P�A� �P�R`<�)�qE|��+,���x�Slބ�$/�uln3z��@��.�#SH�+"'�iv-J�F ��?��JO��5�V6�~0�pM�����z�	[���(r9���j2��ghZ}&$]<�5��LETO:�K���N'�8���*�������J�"�}pZw9��ȋ�ɯ��q�V0�A���3��~�_�3h�hh�+�\��iģ�sr��"���:�y�>V<�	���� �A�����bD�xG���c��
���M$���@�^լ�U�-���Z��0����4,�W�|Z�r��;~@����ߨ}�	$�k�Q�O��X�X�������Mt�@�ǝ_�"]D�H�#t�q�!N:p$�̍��]�؄$p�_Լ�J���JL�pt
�z�R~ø�ǂ�Ow�C�vlO���{�IR��S28���I��9�4˪���o-��zI�F�'�vɝ�*�D┤��zl$��������սF�Fv��T^S�{�3��^R�߆`�<�641��������n�U"7�{��
"��	��5�xDM�cl�"�x��֠/L�I!P	I����)+���O�3
����t�~=�ǰA��`���I��r����Y�35���b�#�,��f+>z�lt-�?@Ȯ���~i����C_��m=� 5jѲ�&��+>��Sh��{��)a�e&!��B����Xt����ճ��$n�@�'�iߙ��X�J��.�(<&��׷J(|��N�Ik�?Y�y��R�VI\H@(2n��^5���$`����m�!�I�["�'�o�C�a�r�ܫy��),�|��LȈy_�
���~hv�K �~�H#)��fS�����J�;��Ϗ	aZ6������z)_ܱ��u�ӿ_�{����3��죂������2u^����w�1Y}�$�Iݹ�}�9�GZ�xp�#��?l�F���h� 
=q�S�s>t�}�lHT*I��r�D៰�A�Ρ��w�F��Jk��� T>�NNA 7�|$�Q�h�&����ǈS��X�ٍ�����C�Ƽ�rN�qr��f�S��z���bl�DC�oxn������fZ�#8qb�ٔ�I<y�\����tb��{=_�+)G�{r�hUy���t<J�����ֵ�tfU6s$M���� �ͪD�{��G[��#�M]��:ȹ?�5�;�P��XZ��u���*qF��[�bV��+�GN��H��X��FT$f�~�hL�p�׀��JY�K*��,�����6!Y�KT@���?���~9�yN���C��nAh��L�����mև�3@�fn�Pb$Kpp��!��M�d4&��<U}D՗h]8��2��]%m�C�?�&�jC06��S��S76�����i��*����I���-����E�@e5fk�����"N�AeZ�>ѕ[�?��Np*����ǋ��c>�ј�TP����Iz�r��Q���ѵ�1`������#��L
ƪc ^�OM&��9e��,yC�}v,��i�����;©}���ii+Dh4�c5/%���3�A"��8�G�KYq"�J�SFD���y3-y�eU�gui�	��8�z���Ag�{X�9�`t�!B���*L~�|e�� gޚ k�o��=nΤQfn���i���GR�L�U�d��}p�%��~�����w����>/�aVL��X�4j
�qv/j����_f��p�k�K���x�A�{$?���m�����S����r�^�ID�v�Fd J�*���V&��~@���Pf��2�%���`�Ф��;�o��֘�Hq=`��Hjl]�&�u)�G�J�a,רn��V/|k0��>�1�
t�N:���t�;9ֵ��X�6I_��A��r�/$b��
�\�C��nL*�&͹�]l���p?��Z�>[n�T�G͝S�|s�;�z�������=�r'�B${�ӎco)B��\���:�qʤթ��g�q��q� \��i.��uׯ�Q�0�p�V�i�e-x�8������*���t>ژ�v��甏¸��?�>q�wj�I�h�EX�D�k(� 	jև�-�.�@�����ʍ�9�E�=�^z.��p��-���p�P���W���p2��k�������cY��?:kZ���a���Rl�$�-'N ��n/4�*¤��Y�/	}5��e ����-�ȗ��asiT���.����#�b9�E�L�1'	�_θ�1�	6{�ah_^#8DP|�D�m5��o�z��Mi� �'�ٽ�?n5G��!Xn�-[X��!�3/V�t���ո�|�^'��Q�G��1u���Ab�r_�0:F�y�5���\�0g-ᴧw���3! #�q�0	2F���z
�².#4�n�|��G_�(���C~>C��6�{��#~�x�X�4�����]�!���!(�}�5���Cg�<��cE��7
��N�]9�O?�����m���*��3�z/�j-Q2���ҝ�:�AI��DӦ�&��w#��m�\~Q��c�c���p�_����z�W߽<�ta"K૩5Ӌ�
��T���r7�e��hx	Mk�L3��B�u��rmDȪ���`�@Ӑq͐5���>.�z�`'���O]]�~�p�v����T�.@����G��j�����5�V*����nu����'z�^ao�|�o�}���u�� Z�hC���|Q�FUy�c�;W�5��D���$��K(U�(�} �*�J�NӄD����_�4<����i&<Q�
��[z:͊�x�*(���~e��~�d�mL�%h��l����H�1�آ�F�r���u��n��s�vk!�k�5������~M��O��㹈�fM&��d�[y��nޒd$}�����Km��Q�j�*.�����$�!(	��x�)���'�c'�DI:78jU�U�?��U��IMv�&�q���6�V:y�[�vn L�; ������Lֻ'��1���L�uX���!3$�<�'���lV-~���DF�:�
�>@%�ȏ@͚6u^��Ѐ"�)�16�Ġ~D.J�~4iX��}�j;Q�.�V�ָ��+��S�z���((H�@��*��8�%w���
7[�L�=_[B5�V�Xw��U�E����j��'KE�S�_�kPȡ�S��kz[&��ۧ���R�ѦY(x��֛��r�d'�����|�p�A?a�*���$e�&P�&�}�`N/��iy�ڋ2JWG�z~>�z�+*�"�ő%�[�q����Z#xD��#.	����L1�4@�P&K����,� Zp��{l�������S`��$�,�����,E݁��5�*��.�G�S�!(�b�y_*���z�G���*h�
ԍΒ�N��#�N���׽���؆����;�mĿ������IY�t)i�d���I@(^��^Wkf�,d��V	\ٙ/�!2�DA$ʂ�.���
I(�<����+��ǺjB��9f�]�<v$��'�B��~�#x�"x�5�9��p45{�M喇��2��q6���X��/N�3��l��Fjڈü�\�l����g�`	qĚ��=0�=�ߥ:�xwz(�_�G�Ó#�~� ����혙1���xbK�k�I�(��1�N����K��t%�ָ~@a_�9M��x٧��� �������]*H�Jxq���M�B!�4���k���E�B�����ec<~mr��}���|!`p��� � �����̽9����|n�H���i�Hw���<~�R���oɁ�~y��eh5���l�^#��f¬�bIﰱ��Oj�yn���k�(��b�='?����I��`.Q�}�R/8��3��7� F%��b��d�����5�c��W��l�vDKI�2]��14��gd^����Օ������ar�0�l1��fA�N��j��0�c[�E���ZF� �'��L��ކ��}�Cy�p��R膁�.���c��v>��䉿�[�2��|������;x���˞\G�������-b'����v/G'�.��}|,kO-p���_g��GD�]Ak$8:�4PNb�;n��7?�M�a�"������r	BA��@>�m#-Z�9�ӳS��"`$���1����������(K�A�b��M+��&*�J���i�}#b=�R���߫��P�J��	e���ҩ�m�R.���8����9��������y2�3,����V�*f���7rv2�ǌ�D���D&-����%ϟ_*B�����ƚ֯4L:w�Xi:��xx�"����n��hsՏ�g% )�]�n^�R[,�g17�6��	X���ߊ@��ϊ�硅aql��l�ū�`���F�WZz��Xv}��Š�)���ݬ���	�j�X�\.[c��2�2�ҷ߸�~���|�r�7I✂F�P��}.�|��H{,��1�4>^��ax�\�Վ�)2��fh}=Kj$yc�V�Go
�ʷKhT�ڨ�%�����(���|c%X�e���*�*����c~��%?L��-dM �����l���r��d�Io#>��d]H�1Jy��Gg!Ը-���g-�u�'�)���S[C��_S�����B�M�v�yC=i,,@���,��PXc��v���1�T��(Ǜ�zh��%+��P��sC�0��&����1�V��}������
X���柈Q�d�m�d��֚c�5�j��'�6Y�)2~~�����n�0�ȑGc��@��Xݏ��al�z ĵ��»��6ȣJ,�>�h9�ʪ�|���l���
�GOӭ��r�g��qsk��gK���WZ����e8K���H�D*R�|�C�����sL�+K�
^��%'��_{���܂�Bݮ���;a(�,@��Yg���z]�L�>;��넮P0Hݠ�*���>�Ye��� �\�+mXږ���������ʔ�?��U�� 8�����y��DFL�7n	�]r��5���R���v���S0k_Agp��c��eχ�?�J58]*�b
��7I#�qpth�D�?� ���'|1�7h��K_:�����y��~=��3��>�w���?�)y�R[�^M*s���m%nnE�" ���
�;Yc��[���x�u�iO�f�͢�=s���
�S��Ů=gi�h�;����xC7��Xg�	Z�s���F�!�o�Nvڇz�����_,��3_���ɻ�_^�37��4
��A�W�e��TJ�:b�y�|�ϙ��F=���O"!�6��4��y�y�z�c��&�M�����W�Q=c%62 �]\�'����#��q�
G��ز�͕��BY9d��x�_�O\M�\٤q� ��B`A�͆���UJ��R��Op�z�c���B�.S ��c�I�}��� >����J�;���y���j_�)zh�e��o�KTy�ƍ��fOd��ʚ36}�{���Z'#�xoz>xH'Z�N��e3���gzk�eA�rm7�#����z�2a����	��.��_�i�Ko%TT����Y� �]1�S��,��W&q�m�e>����%�0x�nOꍅy�(@Z�n��o�7Nv��=�'�d)I��[n�?�;�5X�3�_6i����\:��}u{�lf�N��{��3?�����E֬u���lt��T������g�d0�gQl�Ȫ��;4�<��������߹5P���5"]�gCH=�kAZ��Z!)&\��?D盭�;�IE�7fI)�e)Q��]�#R)"��b�������'�ԝW�LZ���x}���7�-�L�条�$Ŵ w>��[�ئS�e����q����sb ���5o��?6`���m��9�m..�1aQ����EҮ����Oi���x��)�k�K�xJ*��2D̫�s֜������]��*�˓��v�r��<�~~�"��/E�m�M�C=����%f�2��u8����=gY�%�b5�[YQƹO
���!���+�o�
��m_+������$��8���p�aEL��[��� �c�7/��u^xD	���?$��P͊��l)�vjм�c8��2�ۄZ�,w��'������9�c�B�G�>����S����дJ��6b�ʹ�}�9Q]��2�ޏw���

Vs��t�N�_��kMɑ�}�Ihkh�60��B?Ѐm��A�ȳ��B-H�v���5��ɜ6�5�F�,�-D<�bX��_�č�ȉ��?�
I�}��Ү�A;���B�"���}>a�¾@l�Cٵ�z��0�e��<9�Q�U������A[9%�h��]�2�Ԭ�weV��"��p�\�����1�N}��	=��k��=[�o���s>�Z��l9,G7q�V*Z[�(RV9QԦ�N�GY(2g����~��om�E:��du���,��U?"���	G���f��4he�t.������N�J�y��*i�5����m��5X��F��������L��M�l�\��;��;_E����:�f��w�y�:^����E�꒴�.�9���Ie�e�B6H�dP�~��'X�te�jiNl�mJ).�Btq <_)1m����D��5��2pT����Bz���l4J����aQ30�c�i��jK:s1��PI��.�A�J�H����i�Z��Ź��Mw�y,R�HjP�$��#e��ǈ�<XL�����ۀA��j
?`~EQ�J�X>��QQ����c���(��-���8>W5�(&``�g�{o]���E��Or�d���wT
:6�+���-��'e7�4���r�1ܝ-F���Y��5�\���3;N՞�FN�I��fm_ю����I<��'J����VzX4�����߄�ڦ�oZ+3�g��BW��hgY��S�R4Lq֛x�y�����t/5:L�0�$$h�v��sI!c�AL93��*��;�Nw�d!{�Ϙ�Z��ѣ|t@$Ѕ~���)HEq�@�c�XoI�M��� [��`Otp���/ʘT2٤ߍf�i�̴P-���r�,�t�F���Z�!TX���ԝ`}B4}lA������b�T�Kkq������=�e����*wu��c�ӓ�^��&�!� ����+6�"#��"�����A-r�d��,��%��Ǘ�0�PR�Bv% �N�U��tt� �2�_a�k�]t���N��~�1�p��q��f�cNE����x�8'DtL�>�/v �1ѻI-'��I�A��g(:��1����2��e߸w\��ި��N@!i'�ki����t*��a�ܻ�FLe�a�h;K��mJ��y՜��Z�7��͚C>���̩��ĳ���S���a	ނY.�%�}hB�̊�r&+���b��ڒl՝(e�X�.wD��j��� <�࿝�T�_ �6��WEaNلM`�k-!�8Ӯr��g\�Ə>�?�iA�}+[Y��FKUf݁�I�A�t�ͭZlwf��թ!�,`5����D�8we9��1+j K���"�c�OY��Ი�z�������}��LX�	m��/'�ς�'�3��B����?���ڹl�{�n�뽝�߲���)��A�x��!�]X�ǩ/�E >�-&�Q�61b�_hl��)`�]'Y�t*���Y ̼���,�������`��e\�g�2�$�ɘ�{����+d[�R��8 \�/m���Q�W���M���2Y2�G&��ڒ��ھ���엣m�Wm�-o��B�OU�m?�5��U!ݑ�z���IdU���	T�=k�F��_�:J���o��~�oIϞ���EN���9����w�A���C�X�8k����x9p�3m�-;�
q$ٕ���rO���?)r��`�tËY6��k ��J��:f^��̡I�H�\��p�N6E�K͟~�������#���ȩ�i�gL������>pڬ���2�綩,7%�h��b�\���[��R�[��%���3V�p��r I�'���+؞V���tv�N�$6)�岣k�ð% 2���&�..��u�P���d
|ί��.�5��'���=�$�����2�=�x��:�KFUb?��a�_��΄�싸Y�1-wO�[�x���JD�)yG��m��"���v[�]��Y��a,��xdoғ�(� ɅeRӽ���<�Y>ժ�h�K`�����R�0*-d��?����]6��׼�dG��?af����>V��&����ɞ���\����tz�Q-	�,�^��|�G��q�R_\���@���n�Q;�.O��D��`���^NS��\d��E�'k~�1wI�d�D�O5w�bI�#���!�Z��^�Ϧbl:��"��^��R�(�| ���p�|�7��zy�Q����^�`�	F�
�al��}6�3���������)6K�R�YVu��x�Q��Z�Cy�.�U�M�:�)��a��Խ-�n@�d��ZS|
�+��X"Gٚ����
��s8Ǧ���]<c�n��	7WU�%T0����� Js�4L-oX��yecdC�c��h�m/���ht�d�<b9,@b�T�7+�m�È�CX���|,�#FZ�����`�W|9�]�\�[���*�.�����ߗ��%�1zm$�z�k�u'x״�QMc"������Uþ럣>IUSU�S����¢&8r������#��pH���UB5��Wi[����y���cS�(y~���5&Nhl�R|����5��p����	U��>��� ����_��K`�𻫖�|�7I;F�; ��3c����"���Y+�����m"Y<@|��������W�1(+��!�ŐHu�*kx^M^�<`��o��W�E���d�V<�#��	�����m�Z X����z.F��O6aB��@��ϸ?; �|/$y9C��=
��q%�--˨��$���l�ލ�� �S}Z�r���<˩Oio$�Q���!n=���̴�n[����H�H	;��	xL�P���"F��u2�Ѵ�f1�=oO/S�� ���@]�ͦ�
��K���p�x�Ϊ�$rP�B�-�0Zvaa~]2Y�NJ���^dG��n�i��;���,�W'�8H�.b��x?�,��R����u,�f95z�i��]�g��J��دط�b7N;��Q�G�U�9M�M�X颿H,����[h����@�|�z���[ �ɫs/��K���M*(	ؾ	�Xi��ܺ��\"jDG�����w�?�f��F����F�&�(~a���-��X�kg�v?�Ϣ�%��{�d���O%\)X��;�J���u�ƹ�j�$.��R��w�ܓ,$�'��z����A���C]��8.Y*�R��ZpH������o{����m4g�}�%�ܬ�p�B�Ǎ�D��w���x�չ�+S�����{kH���__3Wv��P��X4�j1�bv �Շ�9q������]���fy�W&	F9����Cn�e)<ی��j��1�b���8�"��=3#�#3�͵�(��G>ޙڍ ���BΊ�ҡ�S��©����;#���s\Ϲ�Ο�51'iV:qw���-r�m��Ż��P6U(��vj��������:m�v����n�)$�3��B��ಗ�Wq�"���m@�Ҷ9����;{���P1��<�|�;�Lڀ'̙� !��oI����)��g��&�%�6q[7���
K-)*�O懫�B�>-]q�;+u���d˸��EN��W�M�ء[���y��4��Q��b�%GA���5ʉ�H��xh�.�aF%�#'ffq��W��z
��RJ+
u��� E!Q�� �{w���:��tM�X��yM�8�p�%�oR�L�:�(:
y"�t��K��0�i�y���i-��0�<^S�%nU.���K@c�b��䉄�%RM��#�K���F��	�l�]م�����+�b�<y��>��lh-��g>��i�L��:wrC���|(f���h��̨�_7��+�+��oB식i$���yT"q���ۦ�x+fx�������Ǘ�)uY���|Z��w`D]��9&U�U0��e�����9��6DQiߩiB������G8�#��(��Pt��L��=��AڟJ�ySa	����a���5����!y���M�A�.�9�-�3b�eo�Z�椭/9Uu�j�q?�)���:0epAf�,s$�Z[��OR�uw�v�j&9�[i�Utv)i���Z}��ռ���ř��,��䮎���İ^������hw�$��t�ld�Xm������`� �
��p�5��B;z�{7��]�ɛ*�]�;�Nʭfc�Z�)Zȍ`6�:;	y�I�[�VZ�����Ȭ۽*o��^�р�.?�2J���M��GpD�[L� � �6�"g:�}�`5��ݣވ����{�&�V(_9
0���+y�����|��UP��-���j���֜ő��Ok��V<�/ ��O�ûᲦ����LE�l<�)���76���;χ������
<q"T8B�E
�W�Q��s_9�������c�p�Q�t��O�Zp2�&��<}����|u�9��œæf�®�z�?��bD��`���@�#�n�"*�J���m=I����Оoy�.]��Y��-g~��� $eZd�B�v1M%�o�m �1�l�'V"����]-M"�@d���ǭ]]t�S"'/��e�Dc�����5�}��63�o�p wm̯}��Hn��jLJv������YX�#-n`@ׁ�V���.�x�Y_5�)A5j��{D���洛��#���Cw~ʭ�i��]fG�2#F
{͍�A�fE溺����e�O4�M��%"���avۊMZ����?��~�;Dg�RitCb󠻮U�nz2ˊ�Z^�vR{~��R����y14��R�ک��8�k���R��e�d9|���CeB�֘��^����K潬f�i>����ix)��*;-w��40�H�+�3У�?�`&ʾ^�t.�W�t�qA�22po����K5�
��Z�����kly,� ��\m8�_5pC���.��~̟��k�%]�P��5�����9,��8�uH0dz�;��m���M$k���M��M�> ���c�6�*h$�`1Q+%���IVI�'�_���|G?"�����B��x��'�M��u�!/d�Q%a�J�_&���[���x׿3��|�!;ղ'q`���f\
Ѯ"t$O[��[��A�K����y'�	���T�"�u��D��l 6�^n��l��R�{����yBʄ��.2b,��#MVLr���1���s7 H CX ��t���W� �R�]!
I"ϣ*60�����>�2�'��P5� z���7u<�ůN���qm'~�#��.�F[��.=)ڼ�wZ����h�F����"��w�b���0�P�龆�~uq3K���KU�ED�A_�z�Lc���V�|`���ֳILu��2vV�P�,A@I�r�D&��'Δ���j�|�{{�����΀��5z�G���r֌�_$	���;\�7�C<+��G0���e>m���a��W��Y��WhR�X��.k�?���6�!��۠_#�i�M'��������WvC﹢yޜs ��X����C�]@�E��~1ʨ'�@��Vʨ��j��1p^)�yrF�ؓO�|]��P��Z��~���:\_f�F&�����JF!h�IfL�Zk�A�աVf-I��W�F-�]�:�:��w.,�s�;���,�͛-ʌ�]y�h�6:/-|*lt+��C[�T��{sf1���E_���J�O�cX	���D�n�����}�x\)�wԩ�	ɰ�,���Ke+C��	�e������|�i���NS�UQU�t�p�*`���:���L�p�������.�Y罒P	�x�X/͹by��t5��)ޕ���A��h��Fyx���Z5M�H�<���P �_��:�9�![��y��F�Ux�.� a�V��j	����J����$P�}�G��IDM�Dyӗ�xOM��?���ߏ�W��K�#����)���Xh;B)�saI�M��+������M#ioB��D�$�f�ʆ�D�����S����v����z�&@���h���>v�E��� ��E�L�Z�~�6���Mhi�f ���O����g�8�% \�E�Eq�����P�N/�,�rVU ���z�eЩzֵ�Y����v�O�A۠{������޷&��l%�y'�D���^,я��]m������8Š��ьb���-ʏ�8;��2@ԄR����k}����n5iV<�T�r��v����� c�
'�Ȭ3��� }�Z�4B
K_��'����[�'��m��Ħ=n?�R֐|j��᯦Nc9�v�b���-�6�{#9�a���Dh�p;�A�?X����B�
����Dk=e[�bGDv�d�'������g����I\��=�n\�*&�
*�ЈpǾG�G��+�Ϡ�,�R����>�w�R���NI�Kɀ�����^	�Q���f9���ɱi=�$��]L��پ3�U����t�f}+�L�M�dDR&G�3Ѭ��kE���/�0�*�'�����[2x�E��cE�,`�����Cˏ+eKFn���绶M���{����� �G<�3Ճ���oA�Ժ��I{���Pċs��B���� �����` ���#���}�j�]�����@YU��M��6�ݩpl�H}\�n3fvZHdc:�c�f�N8!��8��h��^9�<n&�Ӿ�we�琶��sWzM����
W�R,H��d�  F37
Ot�G��ȯ�\��kۨ������sY��"�9%���-�������Q_p^�8���X(^����7��"�d��l��* �#]�]��\fߛ��)㚱  D�$��1���D�}�	A��(r()�s듻������ic���\�������z�5W�$5!�k�Ÿ���G�:�B'��1F6�'J_�Q�2�V��u�P���Рp��ʋp���
灯�bxz��TP�Ӡ��JY�l�O�C��2"�="�߶u�{�٥{��| r��ޢ׆�[M���S U�{�U6u$�~X���w�f��r`��4�)'=�wX'd�z���i#	�.�XVPʫ�ᯛI��i����w��l��|D/�"�~Ic�o/�����b�s]SW�C�Γ�S��4�D<!2����V�}2�/F��F�֪�87�^ �ʳ%8�B���~��d�B�*�_w÷xd��9>xU����d����Ҷ�����9��'�	�i�U���2e�S&�������jҫ7sx�8#���ce�WZ��f�_�������=2o��{��:v)0��ҏ�q�0c&�;Ӫ����q&�^��	�eA���<Fyl*�ע���lhT�;��2-%(m�7�Rhˠ���D��a��~LJ@1&D2�҂��C�8U��b��s.]z�r\g㲄��E�TeS�6�c�ϞrF��%{(=��y�0c����n�c��t�Ż)�5�6Kt��ͯ��0���n�)?�W�Y<�i8�4��FA>�2�8��S�
V���`�{�6��[����㸫Ao`��|hƾ.p�U�U�|��3��T��o=�8�l��Λ���>?Ȃ��E\(f��B�T����l���7XtS�"�uL���%��Z����R�t���l�i��'��iW�)���jц���׼��<�2�l:�3��)Cq��.`�����~��W"��v��]�M��pֿj��z!Sa���{}{V�k��	C��;:��p�k+�%��]���B�u�[9��Ӑ��9�o�?���aU� ��X�f��H~I$��f����@B��������Vе���]ڿ{�c�����6�����GV?�;Q�?i�DQci��e��ymo��C7".�ϔ�g�k��@��>S�����J%y{ŧ`^q��Rt���V���Dy�ӡ��m��|c�ʤ��lQ�v�oO��A�����u˓��t}CI��3���xYm�;]D���ǿhk� �=�,�_���	����@/Dg,K�L�|��i+e�,� ����hH܁r�4bH�y�L�j�k�u��a�[.�	�7|~�>{I��������[ʹr���7����k>2��[��Q�k��|�a���Z�Ewӣ��T3A�/?-�fe+j�.0��[9琶ޘ�c�oR�Ϊ�>�Ћ`��Ǭ�g7��*�K����ݛI,o��/��䚹�f���o�*���[1D�4�c�k�9��	ʖ�t���X���/�핁qz���rd�+2[Y��_�L�7DoL@Qy��ic�gX�� V�"��G�&;Q$�Zp&�6kzZ
�������3�v�=!@{і�(�����Cw}~�#�ds�"����٫���p���~Gu�\Y�Rޢ��0ɴ������%�۫lOVو�E;:��������D�B��gX0%-3��*'SЀ=��Z�.�g-Zc�������v�gaz�c��E� .k������S�6LC��㣨��.C�*/���&�8�)��Q�v����.�Z9���<�7$%������Z4纜A�8d����"_�P�A;aۙ�C�f�P��v`�\��s�z�]�����`QJb��J��l$����N!O��Nj��i͵� `<���Ua[��M�r�+i�§K,a�!��LPM!��p��Z����(��t>���'�[%:��KL ִ���M�!&Q�
����I}��˖{�V������8r2��`D/�����b�{�v�U�1�����g��*�>�xz>~Q�zH����%�,|X����y>۰��Q��p[y�Ld �v"g'��������-t�s԰��:��Ļ�p��m�9��� 4�Y7�9~��p@��xz�<�s���l���C:��eLPTw����G����?R�� ���۽ݕ�W�ƿ��~�C6��A��t��]U���m�.��:t��<�������d�]eY���%xC��`0���7��|!^�]V��O��ϽV)� `����sFG/]��N<)m^����=���~Ѻ��N��S/=I�����e��"��3hW��f�7?�^~��5�1Z�\$~�D�gJ�#�v"��8@QI�!VFiTige�����'���N�n��D�Ì�$�+#���D���׀4:����i,��i�@�y�#�ǰEz+�Z-~�q��K��ۇ��̀d{��V/�xΔl�)0�P7�BMKv {�y�$ ��uq�%��gV��DgI#��[�s����N���Q}Q
�v�$Me��^�ڡ��*�,���X6N�2S������ 	��2��q���=���K"�m��t�o�����<����n��97pT�?��4�B�F�*V���a�%�v�X~�E_��K�t�y����DӐ� �A�b��,.�J��*���{v��t�@�㍼l2�>�̪�K�C��W�-�����2؃k�E\x�φ�$v��X	��T�yeWbpB^T�'���qL�{~�+v���t��밂$����Zş����[�KjZ
��Q��9pb����%x�<7���OQ �Ņ��D2�-%#IN�f2s9ɖ�B�����N��5�00yڣ�5��RR��z��%?x&K��@�/�\�Vi�61$� >8&�'W����*z!��k���7w�Լ�Qc?Be�����J�O
Po��37+�&��A\���[�tH�D�>�|�>Ӄ,�HK��%��&�h�1��m�k��դ�94%w��c��3::LIB.I����4G�K����+�[㴛��tv�~�:�T�A��5���O8D�V��k���.1c$[含�?��ʼ��u��%���W"�[|��U�6]�Q
�7A��P��_���3�
�䗫����O֛�O�e2�[>&��}X�@鴁�q6HMR?������M\�{�IX�T�D�P:^�$���I]�U�����e
`GJ�*��R�����I�>ckʮ��������f��<����i�SlW�����Xm]�e�k�e�&Kmk�@\�F��'6�L�ǫ����Ǜ�P���kb�.���k�ѩ��)ǥR~
�Z�|VAF`'I��PL�����.D��Vy��6͝���D���w���#�@QY��1�V����c�6C��z��)�*��ݍ�w�z�?qO	�1I�J�
���tq�I�e8(���1�>��	����M̚��?����R�a�d��L�C�leÕj/��U�\���~`L�������YfF��{z��ݜ��
�*�pS��#\8sl�VS��Fʚ�mO�� ���y	JAN��O'�-�1t������ب�|B���s���_ݫ�����,=��P�ר�-N��}<L�K�\���.��<B���0{�*�r��N���q��O8s?A#�`6xz��P	Y��XM�'���@�>��x�����l2�����B��y�8:�� ��6���;�U���0c���;ak@V�<���W���qނ)���#��I@lTg�]���$�=�{{����f���2ҕC��_� *}[B��叏:v.>��tR�mM�[\�)�j��f�B�o3Sw��_�PZue�r�S�k�eY���2�;Ղm;(JH2����jP$���A���"��?�\�pv[��q�4Fr���C)VS����0�&������|@��&[�z/�iP�r���Ws�Q��x�m�� "<��a"?�����\�Ç'�a:���B����4l�M���]R����8���3�b�v����9����嘻G��e� ��4m�^�N�'Zj�CF%��e�։��O�b�U2]�w�w`��}[b���O����������38$oS��	�=��I}���(��A���I&�Df$���E��+�&S����"�"_�ZZ]	�H�m�	i����xE��/d���ʐ� Л�Ch�9����i�}fj{3�����ܜ��1��FM�;5�y�(����Y���-�w�b� ��ԛd�}���_O������ټb��m���|�Ȃ���%\��5�K,�~2���'w��?2d��7Q�
��$�&z7��'2�:���rf^�  �<$��	�C�q�����^0��{H;��m����̓n����VPɪ��׎>��d�) �B*���\J_qUi��J+:�F������"V=���	�0x��@�r�1���]����j �/��d���8��J#֬d�>$���T�*����I����[aP�^�KUc�'�����ê�aZ��ԓ�l�UX՛#״�\*a�_�n��6]�1� ���Ad�O��3�n�1~��F�;3Hwm�?��1Pҳ%����ZL���){�e��)[�Kс�����B����\���K�?JmG�V)�@=����@�#��e��7�4 F7<�Y��*��E<폣��PsCf�P��a!�è�|u�ݒi֯A���r�+B��~���n��8�輣���H�I�̻RL���*�!��8�U��u�/b�.D�·r`Y*ۜ(�ҍV
}p
��UN"����t)1������6I�"(��+�6�^(���L��!����	t��vM�%���3��C`<9�v#�[��wk�wm������V�>����-��W�s�$%B^M`��3ˊ��׏Jh�B��\�|q��1Q2n��Zؑ��0<�
��b�D<��1Iw��hcewf����p����ȑRi��'�`ǅ���(:�U6}ql.���q�B�sn�u�����wuH�U�P�?���Q�>� M�n��k�cy�\@��T^��<Z��ߘz�$��/�����º#�.����<�tZ� PXw{�_���-P�mϲ�u�e �.-!��ə������\v@�l����yu�B)4V�j��N�|@�iϯ>�t�.��u-k��J%w�������\]��֜��B����d+���F����_�I��5����iu<�t7� x�	~0���]p�hF��ڄJ)٬�s]M^����s�{�����90{��\���	��bۋ��C+v�&�Cb_$��])�E2uK��U�q���yn��mW�"�������?y�d��0O��u��y�|v�	Pϙz��@C��n
*�>ݟ���Ms�S�O��~I�d��S�����d�D��9Ƒ�b�U>��`#��+Xt�«�΅(|�O(���1��9�����m��R	g��5�[i���t4m�Q(��pP>x�L�ⅼ��
|'�����I�X�`�E��`�Pa��h(�~�������R͠�������Tx?�<|B�֔!��mC� �ƫ�>��ҧ�gG�Ě�L#�u�*:Q��F����NX����_L��.!�L�:��X5�T�h+��F�m�1Q�=�y��n����%����U��N��վ��wZ4MMK�D9]8����5��]a�{��X���^���x~�2��}��*�]��OA�vE<��A������t�l��qCM��_����M%�e�GAz�X�c���t�0��XDT���Ac�;&T.���~�&�ð��#��G�9`�\7�!���'..4ױ�X�eX?�� �B0��ʞ�դ��PѓF/C�z{����1�@��zJ:�a��ShV�=d5"�r�� p�˶���R7�Sb���>0�-dy�\ŊuKɢ�s�B��Wn��#��0�ہ�(�1�&�+X3�s�2N��	� �����ļ}��il_���� � �e��m��"=!�<a]ǹd����]5>����G1\����HL���M��g� ���D��,�N8�8�mK@K~��:@���1L��:��=	�R&�O�涪J=�2�qy�<�f��=��O"��R�ܖ����̢*_q��Eo?�-	5��PH���w�X���V9߲�'n}��bq�U`�k��sbI�/x�S��tz���w�O����(�۪6Ï*���!\ؑs�����=��#P��Ў��b�hʝ��z 	��;-g�J�&��^D���!�����`�[E���O�YKuo�����g)�`G��_?���&�G�}����E�d�!}z� �V44�oJ-����^g$�ڳ#�
�/x��n,@��A)�
Gt�$���#�>=��.���I�8rc�K�c��s�*
3,P�f��p�V�R@�8Xq�iM^O[@��9�{��m��󶇇��c�Rݟ^��O:���F{�NCVG�}b�+��8���y_w��x��:Рv H�vm.�� ���l����t����Dڶ-����hPp)d~5����7:�7;Y�,	L0�D�;A�,��e���T��%�2#�>�5V���ϱ:�qx�6��L�I����E�ֆ˳lpk�Gо�ʚp�ǧT6�?*0v�MI���_-��q�8Q�n���[�E�a�rÎ��ƀ4�U~���P8�'�w�h�z%�iXM�2h��h�&M�5�R�֛r$�ϫwg�گe����u�폾��o.�f�J�u���R}ּ|<w�Ԛ@��#e+N
JY/�R�·���h7�E��ȧa�����܄K]m�O��':Ꮺ��ߠ�i=8p�\��Y�dC�k����!�l5�P�>�,���
j��S�k�r^Jf��I��^�&�m�?k���8I���*t@�K�5��=�꧆-��fR�C�,<��u�ᅖ�0�neI����C䵐�ߓ���.�ω�BO���OZ�ͼ��UU��e/?Y�?τ�����J�\wSay+	�E������$�r�~%��}�,f�H���,�&XŴ��+N2E59{j2o��n�b ��>��>�>xԊ���g9�ձf�#ݿё���߻�
�����]Cr")�Ϯ���2FB<+�Uc��*gL�T�#k�zٸ6�n,ت8M�U�Yoomz�V��~:��\��kd�~�1��ʸ��{C�ר�K{�mQ��-�8O��#�+*�Ʒ�<�x�ax,����K�$�]9S� ��W:ৰ���}���z�1����O~����=��ӏ���L9��5B#�D�~��{�' |�)���AE�X7����hv����W�� �9ɿ_�cD]ã�\�s�r�T����?���(��L4���.)��7���n;�˾v���w�5��o�N�)p���F�(���;;�kC[�Dfܶ?d����7h��Х������nW�� +��GeɁ�Y�d�;������~�.�?*�������cDo8�`_'���$�ȣ����WOGz�\��l����Y��f#���N�)&OE^���e�!`i��h�Ux�1�ܠ=W󮚔��� �7�s�M�Umc�1g�'oT�ઍ�-c�����(�����Ԭ��Ǜ}��,��>��l6�%�tL��&kh ��WFK}�y�pc(Ά��n��cQƶ���ؕ&�QQ��wi���'
��7�<5�>0QW?T����IS6�����t�U<A4ë9�ѝ�X�UzFffSl|4�ܱk6�����R�%{��1Nז�t�3�S�X�x8�tI��;�lL#.1릍$�CS�Y����4����6`k׈�=�<�˽�O��g�2������H4�:��uJ͝$�m��~���G�ep��������9�hRx5�3�q���p6�O�-��cH�W?P��Y1�n�<�Rb6Z��C�$e��fĢ��Ega�c�臾C�'N� ݙ,po����A���@�S"Iu�A�M�;V���Ɋ=,'Z�(����?�F��f�Pe�ZhO�t<����ƭ��q���)$nݕ+l��x'Ա"zC�j�>V�4,��}�H���;wauҮ��5ݟj�%�����5G��0�Ъ���%��	���.�5������(2���-h^:��w�4h���<[����N�k���*��&�QV�u63�,/ǽk�$����Э���􃦛V��}���4�׷C���\M췦ʎ��k����xt�9���{��9'}����y&����Է��c��Njj�Od̀�<�܋9xbٜ��1�*5�1���t2��$vtE�^8�CW�TB�=�Ջ�G�Y �eVahK7��@�����'�����/���������\3mD�
������,'����v9�_,߿P�S�i������ҨhUL�vDU.
J�������.���t�s����@#�$˨�%+�}��)yעH�M�@�V���P��`l<��^�u-b\B	��+��
�T,����j7L��ʩ�+&�]�ܝ��p}�;Z�D�YBn,��!ތ��#;ʤ�f������q�QKR\�!��.����������)'LǓ��x=fG���3Ղ�`�_��}x���A����g��1��hp�S�[͚:���"F�h&R���K�-m!���s����Ô$]��8Q�51����/@k�@�x?<��HI�;��L�%Z����/����}�;�~�GUc[�Qbm�ڹTP�/����Ԁ�%�y���ߤ0�+���F�ìG��Xr���f���|���~Z���|�������##�͢#^#�M�����ڢ�c�h��o��"�����5h�A�#�	�=��\���������§,F���ur/MU��h^��9.�&�6d����nF^LTK��nOq����81�
��3Hb,G��@�GL�üθ�+��w������I 2!ؙ�݉�4~n��r�{?'�.!���_��x��x(��FM����E�Վ40�ke�l�eT��g�2�5��2~�<��ۉ�6Je�}�^�ֵV���z�<��&(��i����V�]4��&H\��a7��W���5让<��DD���6��9=7��NФK`���޹+���OҌ,S,�l�G��@���X���՟�h��PS��Ե����Ӂ��+l8&��ە��';*��d��b���<_44mCÈ�<8^$���j���-��<�����-
�N�v`���%hb?�¬����{�z�f�d� ��z�,��[���	@�bT�b�6s���:a�(ѺL*HJ��/Rd�|h����B�A�)���y��ӮɰG52^��lՌ����Mgќm�Ǿ��R��<r� �ܪW��ԭ@n[Ze8P����U(�Cjo������6�L�~��	'��h�����D�����	BPC��z�cx�H����Ř��w=4��3lBMl�c�`e�~�X�ӑ>����m[��]dj�����P��֞���Lv�UyK-]��ڢ�N���P�1�����f���B�J��7T=0��J�ĵ�#�Mх�1W�>���ᘊ3ʇC=���L>W�n�0�3?t��WH��r�9ߑ-e�[�fs����[d�է�w�)�Z��U���$�0������w<D4���I� ֙��5/UԒ�b����!E��e�E2s�P��+YqP���ɜu6�Y���Tb���E�:�K�Q�
4$B�H���Q��3�6��@r�u�B每���}�\�v����~�v�@�⌿�����G�b-J�04���L60{TLeMO���bcM�$��\�#P{tݧ#�ɪ���BA�YP4�ۑ�[7b����7�J��w�7P�1�-/��� }����P��ю��m��{ZZd&9F�$�Z�t�pgA�id@82��%��!wZe��q��� ��^�΂Ah�(o�����gU�~���&�N�L�������TΠ>�j`�൐
1�v�[��}�C�0�5>�����*}a;m���^<X����eG��Ӹɿ(K) ��ǡ�fw�ˬ����ƫ��?�o�����VH�#fk�b	����|�2{�j�{ �q��Y���	�v�w)�����e���^��]�F�����^gIVF�U��"/bKq ɹ��(�l�C�.R��7�Ă�Y����)Kt��`��i �58~[��.�f�^�(0d+��{~:��R
��K>��J,Q��.����P��ש cGD�H@i�u��a��	&�2�<�MC��ߥ<C0�q}�-86�A\O/��Q�'ܹ�E��Պv��t�P
�VA�c'���o^�l8e�eէ�c^���͌�,ԫU�c�%g��n;ÄHE��$!^��}�њ���Tn���"VT��M��Gg�z����Ɠ�H̍B�qLж���#JA~$T8�M�^b"v����|P�Z�&���"���	)L2p�)���R~Ə���"�@U��Q����N�����B-��YQ]�����؈�'gs���$&��)���t8Y�
DlY \�m�큉�?��^V�NlR�)|l^��Ǳ��m=H�<�bn�rz�;HS��&�F�4\rV_�;RR�V~�������������@�X��b:&��;h�c�|�����E��-ZS�j=�aM����l�� ��V�3�F��޵��#T�3����c����.}��(�2�kP����o"+���Sj��T~..�m�{�O����s���vXi��oi�ʕ�V�S�}א��VO��>.�.W ^ M�_��¼��ǀ�O�/$��M�;���Ό_7o��$\4� 7����5uÃfP$܌4MI;�����i��6kZ���Y����쟃&��iԧ�`9�����$�<Z:Q��r`���H	�3"�UQ%c;�w�O�g�mӱ��mA#��Mc�X�M`�&V(��cp�S*����IEr-1��):�/�Rɛlr�W�$C8��R\�l���qf�lG�daj���C��� IQV��
�����Ü��r�4j�B(� ��"0eQ2wz�3������.5��֢XO{m���-����M���L���5�G���kz�M��� ����f�f�'��j��
��	�t�R�%�Q �� u�Ϙ�����!dI ����ɲ��K%c�F�8Z.o�
��߫�˃���0���%.W�w' #4�@�z&yjļQ��g
1l�?$����O�P�z�>�b�孍�! �@��o8��㝏2N�H<y	�H.A�♪��Ĳ������Ͱ��.������6�QA��=i��
�f�o��;��+ffyĥ���:/��6��w�[���D��j���fg#����W���e)E���a?�o��7�do�Q�W�n?�۲�e�����"3��$�DL-B�����_�	�ؚ3�3�ི�Q�:�(���4wa5	�Y���2�} &ۗ�'W>����@3k߆c����O+i�X�-)�%}�����0dG�{�D���Vi������'2��0�`*Q�y����b����vnه���$����Is�[�+a,���a�t߃pu^���4����F$_��ypW��tG;O�yW�n3�&�Ī�xs�A�;��N����̥z�ۮ��,�^Y�Ť{q��d.�����!�2�
ӊ87�=�An��k!�� *(��u�!rr(�f�w�y�x�p͠�(��at�)��	�f��N#a�����uc��%�g�r`��4,���~;�(W)�lH�6����e�5��gS���{t�RhU(��ܨ�akX���wʒ�-@�����(���UG9|�V�Y�L{ͭ��]��&Q^�1�|&M���8鉉���{�j��H`�]q�+'Y���|�g/�r��K���d�pׄ�t��9�{-������>�rN�gy�[q�,O�������?(�]>d�8|/��}��%�s~uTN�8�wD���__SU=12uA�O�����c��zD�p:PPd�s��aɋ������N:L�$�6Ю��-Zt�;kB�r���S�5Ab�8���yNC߃#���d�0\�*��G����}��~5�k.�A�DI��Z�~<w��J��I�| u��u��d$�ޛ�ňԽO�gM2lʻ+إ�Ô#�63q�R/�z���ǂ�OeHLW2��)�!�c����74Wk�����Z-2)�&���r,SA���ր���f�JgF������-��ՠ�xTdL3���=[?޻�A!��֥22Vm���c�� M��\Gj����l������<v�x��
sP��(&o�N��Y���`-�����d%����!�5���د��a�s�==@��� n��!���u��/uRLp
�̨TJ��0�?���~��X`Y�yR[[f �B��=}��i��$�V�Ze&���a���!��	��]���mP�հ���F��n������:=�8���4��}6ȆX����M�3W�S�e|�N�/�9ꋙ�JG� ��%_)7q�R�%Ik����C;Y�rc�x�u�_QpL����iB����+�tU�B��W���V�qVq�w�euy){=ڍ,�Q;.C���p�B����Z`B�v�	��R�'�|A�����։eCğ�[	���]f����"6�/��١��d�Ⱦ�"���be���� ���ȓ�ʃ��|T�(^���u6a�]޽[ӡ�W����}
��	�ݲ��8�ߎ�i��z|�b�_8\� ���Gr/m���!�b�8)�Ʌ�2����e5E.[b��Uܿ��QAlWn�@�u� l[|xqv��=4�%���_c��y��A��S�C h�*�~K:P�Fq�+&J&QO�q`�.ϸ��跼
i��������JEOLj�0���H0{YPr�'χ�7�:?��W#�l��)���ם�Ӝ�\|;^DݼV�}����-��wMvpݕ�%�A�k�T8F�DO������e�� ��.��v�ET��K����&��:�"���=��0�5����MX��i����.+���.��I	 �Mo�8%�~��C�<Hի��1��JLdkw繈�Cx����:���R4�$�"t��L�����d�p�u��).E��j�J������b���+,Ǟ�\��=�;Wƶ���;#{.1X��)}�f�J�q9��� ���,�Q�dXp�[=�|z�M2ADe�C�@�z���qGF�@�7��{�${6��.d�q����03�Z�xş�9�f;����� ��*��ieT�Md2�ī��F�{8��q�)b��j�$�Z�ͯ��p!6O�0��v���*S��W��+n��`����ĐB{W]+A^\R��rK;L������X�7+�]F�0� �F����a}��E��] ��p�1��b��P�8�"+�=�d�{Df��v�q�,Q}l���2�]O�u�Q���a�dEO�v$K���S6����m�I U�4nm�/<`�"�?d��̡ۿ��;�'[M��#{��Wc)4ІJ����u�f�����`��X��X�y�5�簶�7p% <4\�j��h_��TV.�g+��I4P*\v1v�v.dDd�~��$�l�%�4jy_�X�V?�$R���h0��]X�9-wp`B]���Q����!!*����ߓCb��~4>���F�|��9x<�����c��3�؈�QA��
���V�����
R	�T����Z0�P �v#qg��D�[���F�~W�(Ks( gw�N9G�C���/����!�0IJ�7��! qI�P�!������'n��*��vw*	�	V�����Q�E �6F��4�t��`�:[O�ă�I��.���X0�XHJߴ� y���v�k�7�$����}�IH/���GIǒ�	0��p���}Bp�,�[�e��A/�**��&-�M�`Ah�J��S�2$��89��8��k��@}c+�>r8z�zb��!�����Рv�FJ����݀g�L��t,����)��\�@��jp'Q��cq�u�邙�xZB��"������O�yzv���ה�]���a�_�V���++����bWW7����j�S���h���=�2(R���m�#�iiq_�/�&#�jPY�X��+�=9TZ��jNy�! ؙ�͊��G		N��"yv��?��M�ع�k �j�� I�v�!۩3E��>�H��FǸ	��ӛ:�I<�x"��z��v�Vc8�+H P[g��
Y��7b��ˆ�_�]���5�5�Ǘ���Ż��66P�ʸ.�`و��G,����D�
��\�l�����=��Q�]�4�T�\U�d���i����]U�v���z��x��8Zz��Q�J9��}x/U��qu +W�u���5�f��Z�����ZF�M�����@�b|3��"�[�R�U�n�dW"���J�s��~��������J	d�Z�o�u~�P�����Ҷ�:��������W�u+  �[~9"z��$��<t6ij�՘i'�-o�{����Nר�����A��R�\-\J)0S?��Y����Y�V���>�(A8m%���M ���O�
T2�����3/�����#��	��o]��cj]�ql��^��������թ!���M�i��M�wB{�i��i$�~�	��#�7�ձ܈CѱB���:$���8�E!wj��OѕG`.5��;�%�	��k.Έ�P�:���_�s� ���| �wiE�;;�\�����J��dq;L�za�fhF!�]K�L�#�D���.�%�s� EX����]��S�C��������NV�Ī�2��T�ݠ��߄:"/ ��[>�+COP»��y��l\~C��hU?x��F�>5k@!�%?�Pȑ�`�@w�]�w�F��+�+^@�h���"�m�hv=~�\�i�!.�������w��F��g3�'�p�؈��.1�C�����޷�Yp��c��,l'�ݑ�2�ީ�r�ìc�D����^�J�:$�̈́�;�&�p-�yH����D ?�a9�,��M�J���;糾K>^]E�=>�$6����-OXp���fm̱M
�g3n��c��SP\�8�#5R�$ۆ�5׭�W2FZ�g7IﺂǦ�-qe�#J`����s
��<'�)Fq��\3$�����#Y(���� x���u�;���#�	3ʪ���H]\h���o�k�˅9��N�� ��.����M̚Lj2��BG򨓳}�bDR����6�b�x>��K!d�v�PX��R����6q6	�o��V�1�Dz۵s�[>YU/����y�M7m��уW�ޒDq.�"w�>8�)۰==k�|y�bW�� `0�P��� ��s�*�s9%�cj��C�ʝS�g��;.��^p��'�H�w��l�ct�f�X�:s���V�^s�ϝ6~d��~8r*e}{6|�ص��쉊��ˢk�W6�H�����_+*X ^�f4ڞ<I�W+�}y�݅,V�s��P�����J����Ur���F{�Ȟ����k-��;9�(�< �1JĈ#/�=^&7��/��j��d�Ԟ,:Н�}�R�<��#8����p�\Чg�ִ|���3���� ���:\ ,n"�DQ~
R�ay'5@��U�[�I�y�����B����-VbJ5GV%9���|�k�[�'�t覘�����=1��iG�VL�Z%�")0�>V6��GcI_�G S��Řdʝ��i�"��.��Y0FlSac���MT/&,�t7)3�$ g�!��g�ͳ Ӿ���6l�U:	UvPu;�U�6~����Q�I�h��:l�2�H���a�5B=�uX>q�z��@j@�K��ԍ��\KQ��{���Q���r�	�5�G}�ij�L>��8�O��Z�n���y�
¦Gvb�n�9���M�]f�f�d�Z.�����໙��C�����+j�"X �c��IU,���L�}�ᙿ�ߍ#+��	3�ie��A#-�U|�B+���x�E��C׃���̬n��d����^�3@�ȟ��{�k�1��:�a�3���)r��K���Qb�+q��+}`�E��{j�gw��7뾛�y.~��T�
V�D�N��~��Pӗ���`2��l��b0x��Q��!�㋋ҫݙ�lxeȐ��D�D�썮LhL���Գ��XMjvN�YH�֕�܈����Z��������c�3�=v"�ހq�D�؜M�ꓠ���L�@=��W����%D�@�Rr��Y/m�w�
b=͑9�@�]�����F��u4�u?��ީ�R!����H�U�ІK�k_Z�;�n��<:P����>�ަ2�=����~�B�O���U	.F���ô16��MLXz6W� Tb������m,�v9<����X�H����rN�����g*���̚��NJml)Z/���gR�]V<ޯ��� ��~�������:��k<HFNY~�W�̰�b��}҇��AmU2��g�Wt�@���oҷ�o��F��{F��GUŘ6��F����LH���X|��O&�}"��ԗ�A-MBXy
&1��v]MTx�%��oW/��^�[�'I��f�[~�tJU��[�`%%|:��k�<���5@ x��c�Ά���o?�`��O��#�딓A>oN�I��0�ƺ�	r����0�Tn��^�����ϪwB�U��c�:b��II�������I]&�NxP�q�c6�L{�Am3�=8�P�eppCoTA�b�ڹN���:5�+R�_�f�<����y��(Y��%�z�ͽp;��<�Tfu�$`d�?�����FA|��t�?c�vq��d�)_xð�k��/��:}�4 /�_�����ɨ�������t�"閽Y��y�`a�AQ��x
��V���yI�IIZ��B�zA3���z�0�"��/�v���H6�q�z ZC�f�Y����Y@a� XH����\pt�ǟ-���O̠��]��>�o�2������3�axm�����JR�ˢu^�E1+���|������ȯ�S䢢?8`��f����Pj!S�4��f50=�����m��ʓ�(��;�)�O��^T2-G_���x��x n?d�0*���>] �p�y���?���ተqn,�cwV�S�̒a����e	�#���ll<ok��V����[��\�pB@��d�r���0frh��bMčz�L�G��p^v���W*�/����^��$��9y��[Z.a��f��d��p�H�O]�Ꜫ�_bed�����W|ө6�KA V� �q4 M9}����.�d�-�I�gUt�����ǰ������o�N>bYI1�6�����*���e�L���H�S`AM�d�[����d���8�<�@��^��,�J"B���Vq��V��J-) 'U1JW�N��~]`JL]���oٷF��L>㮃���pd�����I�������n D�g�o8"9����¥�|�r�9b�����Ӡ�A��.�M��7�hp�4��n��[���8҂7٬B�4l(`+ᾆty�����q������Z >�K�4��=!ƐlTX�M�e�T�[VJ$�����t���?>��Jфeȓ9W2p�t���8�� ��ѽd[�K��,e�L���t�B��[ޣ���ܷz�j�5K�Y��H�p�׵	�[�#�Z�3S(���<W�M`?d�bb��
@`���=�w�c�	^�|��k{B�o���4%>�4^�ʘ�gO,E� ��.���1��2
�
}��w	��jQL�&4��~����W���q��S���"��9>U�0���蓓V��S�ȇ�f���K�uº�:1���<�2!��]�yK�Ӕד-�$��z#��8���Z�oS)R��܋o��k� � �b�8�t��38[D��?[=�}/Q̄vP�^y��gT���K�d�����:��~�jهfV��c�Z��@G�B�ȥ$څ�4�V���3�n���ȱ�y�>��h�66kc6K$S��y�W*܉U� ���@����c�V����
o����1#]�������)�fF	��u�:�a�8T,M�[�i��S�sr� �&'Ý�YaAS0
�k�Ux��_���׉R���S$��Qu0�>.	��f«�����ph�<\q�.���ߔ�q�t07��ob��tk�����O� ��`l: �,��ʋ�]lu��b�y�àƪ&˓8�t?l� �
+5W2-9���C�Mff4o�Z^	;"��֐g���� 3�9F�x{�-�ڊ�f�c�_������/���$m�[.c��2���Ux�MXIf���ǃ�¶�0������=m�]�>w��ܼVn�əbe?����|�7��|�����X���(�I^��1��q9!�ߌ2>�Q]˺�+�-O��G ;�Jvd{I8�J����H��wz	��"�c̨͢��V�cg�݌ �����aQ��+!7nE�Q��Ĭ}��ܱV�~6m�е1w�A���{z�m��~�tfg޷�Փ�qڶ&o_U�T72�WA�C0��a��sÖWO�\�N �x[��V�����᝻I���3��cګ@,E�y�zݝS���J�s��y �W��\P�0H�ݕ��#Ar��A�0����~�j��񟃪]�:5~��zp��R���m��Pl���޵�'�+Wl�+�b�����G)��S{E�^����W��	���5N�0;��h��d6ג�����*�&�w�ll/B� ��b��+�|6��E���'���E2��{��$Dx���,�s~
q�y<OJ6<��T��0���aM�:��c��)��kj��컴�ihog ]����X��4�uO_dؾ�=,WĔ�H(:`G���
�W[u�jb�J&V�a�R�����!��%(5Jo�.	��3a�9��2�/v�dk ��<=Ef�.Eb{� L"��~�X�L��3S���sQC�;vS�D��G~L�P#s7F���B�
S�?��}��N�k��ҹ��t�;���z��O:Uk3#����.����ֆ3H=/��%��ȕm?s�����L��2��6���`���[���Aۈ5|��*I�,PȻ�X��8K�3ӳ�H�.*.��U�+�1��~�����AxbY	Ĭ� ��e2v�LS��%@6.T�7�`T<Wef�G��C5��d�G���!~�u�l�d1�t���L�uZ	���vL��CZ���s<����^4$��y�"�?���&f�-ܟ��\�Ѐ�F뫠�'�)���pP��=�\!�����з�Ĳ��F>�oږ��@��o���Qc�_{�buI�_�q�3헜�D~�A��pF�2���/�Ibm�	$~�_����~�/��Mtv���u�G;b�����ؕ�}M��@кN-�l���UpVzD*��'��ݹ�� �j�KB�g~����'���l���;�S�{�>�:�co%�b�Y�:ha�d吃.wWl�r��^�$p��nC	��e)��3�aR4̝�Z}bhvVp�4��^2���A��]ݟ�+O��G��*qm�,�J�1�@`��(��1zRy珞ij����NRࠚ��[��B_����z�Y)��g6�u��k���6�PE�v>���@�8�H�Eaތ� �@i6r�(�_���Gç[��n�v�lSv��mb	��i!\�iؕ3�lto�X�sY_�?�}]P#|�� �����$"��K�M7P!Y��ܸ0�B�\���n�N,ǜ�JPbQy�[�w�[lj���L�nROەHj�ӊ^ �*�������r�zc���-����KRo��龷�:u�D,?�8y��N��!� ��4�������n�>������Q梜;ӣH�ُ�q�W�P�ך�$���H��PǱp{| `�w�Q�$��� �\�!Z����CW(w�_�|�ĈS�F�f��^ �(8�l�<��Ͱ�E;V1)� (��r=�n�ݡY�.Qy�i7�>����pMH�T�x�c�Jw�,I �ôf)�i�^:�b�ٴf�-�cr�87�����i�����Q,"�f�T��]�)�#�(OV�2�z^��N#���݉8zsz	�s$0�b�&D��&]��6ql�Y�l6%�d��'��-!�u���"}���t��S�>V�#�<�)>�)�I�T,#��hu��C�?���{�-3����������"h,�2��I&ch�U�Ylvw��k�ז�� ����M��a |@,18X����`7�#~k���1���E���XA\n ���\�S4�Ы4�P�ﱁ1Y��gJ��S��y�JPyH��`Ds|��1]�Rk�f�$��) 
7明��@���bծ�3SY,5i�� 6 ��"��M�>��GxijB�J��ܦ�����_���^-x����d-�B-��¦�_m��1��	�\=,��z��R�t-���������ڕI�v��t�1�����`8��'��Y��y��0jZۜ\T��|����%�ބ/�aܐ��\�F��ߴ%��V�
y֍�6�urqOΪT`oڪܪ��O�v�����r�ڡ�����$�r�i� �Uͫ�9�jl%ͽ2�M�V-z�ǘ���o��c��� g"Z�W��lQ�]�+U��	�{��pH >#���W����
��F?��0���#�$�#u)TR0�\*`�g[����;�$�F�4��pe���c��޼��A��#����=���hk	[��$~�Ĭ�\��,��������u��[^$���0>���~�!K&�t ��3�R�C0�Yn��zgS~�ebTl�T�Li��?J�>�(g��2g�T���k��ti!�_����j��'�Iua�>�uR�_7kRd�%!�	���0��,���=oz�]03�=��`7�5���zv���)h�3���k�}GM0y�Y��t��e�H-��X�g�'M��ӻ�jZ�}�0]jF������W�M�1Ԭ$'ò�ݔ��C(�aeav�9�&e�qT��~�.J�㛆��\6�h}9��|Oo�wrX�<'54����M�; W�<!�U^��V��=�C.W��=���$r�扚��9�մS����b��M�� ͉��WD�t��B���|�i�B��cM���V`Y̰�3�( ����U��2b 浮? �gz�������m~�w����/�LzLs�>R�$�R<A	��9�^����m�hE�"1�- `�ޭ�5�L1����V��%��i��o���] MO�ԁ����F��jŁ��\|�g>�w�~t7��h2B7,�\h���]���ڪ6�i"r���ak��c���p�&Q�ebV��GKA�E�l�'a���� =��_�=�6��$?�j��Ѝ�V��Y���1��;[��(� ����R�ˌ$�P��D����52 W(�&Y�
Yt���|Qj�SK$��Jo�`�Qa�*KS!Sې���� ش��#]�j9X������T-�s�i4^Vp$�eG�����3>i-%�]���"����U���>Ҕ��$j���!�?o�Y�����.���d�'�n5�-%�<�v����T
�.�j�/?��]���4�j����>h�����d���r�q�ѧ��\��,w����`#�4�j;f�-��q��ĳ��W��i��|cQl�,l���n��D͒%����,���w,8'ALzS��pJYկ�����g(V�>���L8~��Y�O��)�[���=��[Q�"����C>
߄E;��>�\���Y�0���\1���͹B�l�+	�V�����E)����.K�%�**c�^̲c�˱�e	�q�����X6G�����;�����y��r;/+tt���^���^��ú��&"��DWi�S8y�B<B��v͒�yl�zɎ�~��@L~e�ϛ�Y NTG�3]}Q̚ar^hL��.Z֒�]Yb#f�r>��� �.�\���P�Uqz�j��/2��QƜ����SL��-Wt�����:���i��X�֟k4ܬ�
i�n���f��`���5���L�	������j���>�<������J�b�y[����{��Re�&�^f���,|d�V,��	+�*��8���KP����+��r�N%�9C�]�ty��;���}�%�-HkABl5�3�J������#���`���y��nS���b�#D���Yz`��()�}���?;n�Y��D|D��\�G�Z��_�i�\�;ï�
���ը��a
G������p�������Y����)ޯ%ؽ��1x��Z��p}(��	��kL���C�B��W�sy䦇�d�G�O�E΍aWI%�ty���a�z΋�����/8	��ѬT�I��t��}b������,T13v��a�b��U�]��H3�%��%�������v�L���?����Ɋ��M����Ι�Ʈ�a��c=�0cfA�K)O��i�r���L;�&&k����J;�ℌ�F L����h� y�5ԩH4�?���Ē�����w?B�((`�����v��6��϶�z�(�Ny����	Q���_����ر���G%b2���}Kf�q6_̥��I��j-����A�7���aw�8�s=��k�i��[�(MEI��6��)�xgu�D���I�G{[�[� �#`��R^�����N
��]�8K83���?�e�Jc�9.�BRcf|3it��ijPRB���pY,�
�#��8[��7���N�jS��t�`�B����m�?n�J͇Vu���T歁�u�.$Os�҅9۶)�ǟ�{�v�/�`�e�>@���{Ⲱ7�����,�5�_Xu�]�Z����|�cv$�@�o`%M��U��Բ��
7��j�3�C~Ij{��rۛ4����1I���E��wZ�c*��Ș�~M�ѐ��<�:{�1�Ͻ�{Kġ&$�Q�������[����6eu�b9;�R�&��T���ga����r�����aI5��ւy�ѧ���/��6�v�"�!.a_+�n�{������iقy �c�nNo��#[�a�	�W��q�ӎe��)z��ё{�	M�����S^�y-�:�"T�<���:Hƈ{]�H���Ў�"��D>��mA�M�L-�T���[`��������O��.fJ�.|`��}z�5��'Յ^��l�d�:��+*����Ke��Z�R"�����7�zW�j��D�Ȅ8���V��،��V�c6�\B+Oe��ݺ��2se��4��{眐���7VVAY!L�O�+�ֹ�&~~Z��K�:�I.?)�ut$��6��.���xkN�A����sj�.��\tj6��MN���_�]S�U�r@�uy+5��}�v�R̠ٶLǗ�)���0@��*E�E�� ��"��
�~S���Ve��=�h�����$�JԎl�a@�h�>"ӕ�b����jOXZ+aܭ���S�p��^oM����~?��<��'�����%�YT*n	�uԥdE�Z�����W
���^m��<������Q�l0P�F�I>,�>�L5�(#��݀��t�̙�v��Za��.|���ˍ�]�ڍZ��5���o)F�m8zh�a&�*����j���).�I�1>�L��
؄��B�']KA��u��렆ɛSr��1���~�IK*����V��B�3�y�"�h��>{yg#o����<y,������jJ��o��;3�>X�+3�34Am6ތ�6u!܆V��V�ۑ��գ�D����n"���l����猷O3s�^�O~�O�w?%ނ;2���'�$C<w���-p���#-��e��X_RG4��N[�(�LR�@Ԅ���t��~��ﳸ�v����.ܴ��nmV )��'�}Fr ��)�S
.:y�92~�MϪ+v��e�iĉ���.XH�1o,�
CC[^����E�!��7H�چu���C����>�h�0"$"��]��lѪ��,l�Ԓ:_��P�cx�����iZR�,^F$}>�y=�@mg�Ί����e~���鰴)h¤�98v���>�V�DT�$?���̦��,Bg�)�$r;���TzJH�v��i���I«�l\P�4����!���4�qW�=��7�p�����؛�����}/Zѧ��U��"��JO�kU����}o\���U��9�y$�d �4
�B$���=�S}�J�GE�d4�5��{C�=>o���h�d�N8�zu� ��;�QԼxP.�V��Edm<!P�Wng��`
���J�w�@��#	nz�7��hot%��B@�,D��ԳA���^f,YL}2d�����,�'��?�ܐ��YMP$~�:��Z!#K����8�F�Z����D�
�FJ
��S���j�U=ӌXg_�m/6.��^�|3��?ߥx[tb�m�_�F(D��//�B��TS)�҅�d7�zk���ӳ٫T~j��~��g�ĕ)N��â�H^,���]�"Y�ъt�W?F}+4����1 ��\��Ia�H(��}��I��S#U���z]��f�s]Ra�.^9Î�E�����,Tg�d����Viv�yt]�)M�36������d�~f+X#rMu�Ž��ڿ!4��26���֗=���鿄�R�N�=e����%@b��'F�uG�.�I������r�B�W���.�����~�����#M{6���SKT}}C�v�N�VGL��d�����Bpf�K����V���j��օ����˂"HzҜm���yy�A���^E�D�5��(��d��|�V��faE3��HE_r2���^�m�����%:(�˔���s�M1���C#T�bL��?1�y�����F�\��eGP�����<����W�ƍ깔�>��K�>�����Vo�Ƒb��T����ڗe5�6X1��R�LL7�9B���rjU*<�!w���
:�
D��E�g�[ｋ|<� ?��h,fֳ�m����z&����l.
0�ٴ�~�J��P>�.4L�7(���Z�0�_��3\��G �fTsq��e2�-L�gwZH@����R�tS9�����Xa�ZЕߒ�&��� ��G����$2j2��J�s��/�ꏟgt�̐���VU[s�B���z�Gk+ؓo�7��I�ءM��-{N����MׯP������<�R��7w��@���l�5����A�!��9V����ĵ���vk���JkG�iRP�D�+QzIk���N�=�
�����(��zj�����9Y�B��f��*T��$�Z�Ǚ2[�N	�t���@_:.�����G9���6V%�{���	�A	����uU"x���3ܕT������"�V'gUQ<H��x���t����9l�i�n^'x��w9@���F��>���ѷ��k["s�8�}�Y'I^���C/�[@��RV���pg<!�'�T�Y�.z�%�� @1ӷI��͆`�OϹ��f�����e��f�~�F׫�/a�_�x�(��>z��Ż��kNjT%��w��m���C��>[T�2�P�V���7�q	����ҁlڛ(��Q�{EH~���ݼț�Z��I��<�G˖1D�=�#{7Rv!}H:�m.:�~\Uy>�7�p�K1�f�-ǈ���Vm/WX�/�B�s��U�\�����o>�j0�T�qer�z>�4�p��A`Hi8��~��6k�X>q�tLG�Ŗ�e�!b��������{��}��h�[�'�m���NT�ui�aZ��up�lG=$<1�r��ߦ39i@�&rʋ��6��~��$��.@�}�����Lb���a'�Ym\p0��{äjZ�{�Y+|�YvM�4�VMjN���`��d��nL>2�mz�Be�Ǭ�L�wW\�P!�Ñ�k0}4�P𾯭x��"���r2���W+��L���!��?&*�,h�q@b�4�$�غ�:P�:����8-lZ���w?M�ܟ915�ң���U̩!Q0{{�(�����@��/:��a�������P�5��bg���L���~R�j�� �Y`�P�g�/���rVH���{�be;͔o��a����x8m����3��wT�����neM�d�ۘ��^[��w�}ppMv��N��]�{]�1hyV>��'�p씬8L+��2s���G�
|s��X���V�${D�[ȅ�'.�+J�P�3��HM����+�wk�u.��muJ#�QK@���0U�	0L����
��3}�?��]�;��8֕M�6 �gm&e����_�z�1s�h0�Bt�y��C��z�Of(��Ì��r��t�2�-�-�}��B&R�#�U�N�90�(�i١Z��9{��T�љko�G�W�#=���p��~��	�����;"�%�T��`���;4u�� ~H��ڮ���*ħ|��=I�IT� �WpW��V���#ѡ��t��������y�r!����Wyp�|AF1�Ut��Fڧ�4*�oz�A~�����ծ�ձ�R'���"A,R��{��]�*� �L�t�\Q��-X%C��P}�ե�{VV����F��\�X"ƣ��.#hUD&�4͊XI6!=��^��i�e���qg&�n�:�	��N�W#�j���i\��Ff��뀍�`Z�tK�k�ޭ��6"��Z���o��N�ZH}�(f�v���ZV�Ně'�<}��Z5�P)��r��,���$�MOF_�m��������P��6�!� ;�\.>�U5�$j"�YM�9��") R��B�}��R�)^�r7�\���H��M�i�ר�4�q�-�8���@�5�/�q"����:��T*TK;9{^���ޱ̌�)6� m-�z��IV��G��ɪ�����	���$�ể��!wBi�M5� ��g�T����5��������0�ԃz��q9���J����5�c`/����)�:��^�p:8�֐k�]�Y���@~&�ُH�f[�uCB8��>���s�>�;\mSH�П�i�a�aِ�p���������3��Õ*L%l$O�N���߶u8��N^�^�j_nT�c�z�u�y�����=��ȆF�ü.Xv�9���沏z�j�,�� ?�t�<�i����>�y�>Z��ۓ���Ŕ-!h[�,��0+����w�ocI��!T�aS0�LE�`��	�N6�ѩe��R�7�&��R����=a�H�wו�?a�2?d����dS:�l&�j(*��ά�eo莸���uB������=X:k[�N�rMu����tbb��qQ����t#���*��4�~g�8�u$��!�ZAiқ�^�T0�Ei�o{؛ܢ���JHbF���+Uo~����hvȬ8�̋�'�ݑ �9 l��'�?�{�s�}��h�V��|���<؍*�_sxk�ݹ�$3��Z3�ݢ&�R>	�ʻc?�٤�� -i/�AQ�ӵ�V�bW�>a���i�o�3V<��Z�ց�Uܒ��JJ�j�*��QS�Vw� ��7;s��w��1������=�a"0��E��c�sÑ��s�^ۯ�x��?����dL�:(��Z5^>��" �����?�z[����H����J '>)odlP��4c��Q~f 0��n�iI�B��2��P��?�y����K�L��2�/�q3���Z+G�ԛ,���d�,�-�۝��`��	Mr*�%>�BϽ��T���
w���!5G�8T.����nH?���j��8 ����D�}��G�O�29_����w���������~{���*.����L�����|�"�C�8�U#h�W9�h��P��Z�,�����ͦ!�6Ώ@�F���I |�V*���	ƃ�F���#e��_)��=�������L��h�n9g~(M���r����yu��j�~�=������,��NK�㥃��E�~1�1Q5`e!�=�ͷ���Sof�Q�T�#�0��,v�n��J� �V^c�٥0����	�I�L�
����0���!2�\Q�\Ϲ����E�ݜ;H�������)J�f�N~*8����N��.,��@���oh�sAJQ��l�1��/�`~�9��Ȁ��em��=��G��B���c[o��OG�DХꜺ�Rǥ�#iI&	�B�|1#���V�Vaz�r��S��?�GyF���YeU����|��.mW|�,)� {o���Jr��o��4y2+�d�����o)}@���Lpk�T��H��}������h �1Lm��?�q4�Ep6�n5{C�F��>?��M�T}�AH��̀;{>%b��k��5'h:�O����ؒ�<S�U��{"�o#l��j/M+Ww��9@�aF�U&�ߩL�Y��Wl�bBS����aP��J"�@c�z8{�兝�̸����%F�hR���Ί���'H�[�})X�s���9�>�/�^^͟�3���R��q1�#�o�,n��uH�~׶�z��T�
��]��CG�����A����~Eg(_FWB��7�2}�rPQ�|��iw�{|��x�o��q�my?r���c�ʪ���@}�ս�l����T�z��I���T�y�|�HO�ݬT
��Y�
I^^T�w�[����R,͝�)�*ć�E/\7��T�SKU���W?]1��e��ΥY��H;+jg3��8]��;IU{!�CZ�2~|)��,�F�
�)�.NԆ��t�-%*���"��k�K5���k|�� a�'<5M%.�؉?	��1�݈�Ì-�İ"�4ߠ	"��-t�k\}�?��Иp����p>�e�8�l�dϵw�ъ��ܩA!����^ ��S��ߜ���vG�L�|П�;�DK��AV��|{.Z�h�~<�M���x$���+O�<��\ƫ��TLU��e6Op�����K�D��n�	�06 g̛+sCD��CRS� ��j0�s�,y^_P��G WJ=�jL�	�ͮ��=���*���R�p֤��0�.'ןk�$r����&[Իa�q��t�.n�}A�A7�r�y	ss��8���#�}��jB��4;����ԝ��O�K�N�(�!�6�Rg���� C�����)�5�:n=$���|��k)�Iz��&Y������h�Ȧ���Ce�n=l�8��!�>�� �>�l�[Մlw<�ɯ˭��L�j���5oa��n������(�`R�� ��K�(�R?_�m�|;�����=���J}@P���3`�2����L����ӣ0�yV�DjjC,>6!(L����&[�$��'�w�<j��!`��U�[(�RX67'�*��Pެ���<TK�\ u1pe�?jV�xgs��˿f�1,{ּcsJV��Q������`;��S�@���8SKN�RlZ�w���O��l�	h�hū�&�����6ʈk;�V�������Ӟ�>�Po��kc���0����#�'����h�E+�����zЪ]�CG9��W1�^����^	���0mp�\K)�as��f��a^l_���_9�	Ű�����/"D�ZY�vB����>.7!�X��,�?�*?�n�37hz$�E�{��m����ĳIL}��BVEw=�1Qj�0Z�	�j�qC��,W�w���7V��L:ۈ��|X�R�jc<�h�r����z����:!چ,9F�Ȣ����ڒ@�yez�K��e�l�j�;{�%�%�4��l�2� j��CY��i�x���Z�]��0%Ļy�AM\�YW��2��x��`v��Z�t�5����ߑ���w�	(6�v�k3G�dQ0K�u��hR*��&���|����%�3�ר}^��Rx!�߈ä�Hz��������ho�t�z��YTb��([�>=��7wX�s�k�ڿj��5��~g�m������r0!�nl�}ş.��������ic��54Ќ}$Z)���� �p��L�_<V�}եS6B�����~,���R���vv��xNPǖ�Y���H�	�S!��ޜ�h8�	�fʕXE����W�����Sɦ��Z=�ב#��v~���@�?�.hv>c�;{�xښ<Q�	��{�Y;U;�p!O'M5��Q�F�[G���oC�D�.V��e(܀>u"o�{��!�Ѭ�����b�[����2�ݛ\��( H ����?�)��b�}��T��Q��3��J�a�m�����!�`�>����=�*�{�����|��vI.)C���l��)�[�9UJ�⯏$�Q��s0�(�����H�1�Oa</ P���guI�j�O5�����l������j`� 22H`ʭ�dp�����=���� oi�ٚ`P�ă."����8�*���;�쨍`��R�����(�x�� e��k�%;"�a'��v�8s�&�S6Z�Dp�J@*��+Oȵ��7��:���E�&��dN�{�1�Z��2pm^t��Ӗ������֦��XJi	����9�eǍUC�v��е���i��䲻�<�n�"�X��@B����]<��H��ª!I�� `�iC��3o�+��{W�7su�Q��^hdf�r��sL
�t�v\5%�t�������\#;@��J�P�e�p���i�����a��,�~�CIpW��#�؈V�c8@�o}_%��n�6��z��mBW_���rP��)�Wm`z�̯R�؂���>j��a-��Zk��#"��PɌt�{|X�Jн���q���\]���{r]�{�@�>!��5�7���)[�)���5$[2�m,�M��w�P��.����xB<r���R|�Rlq?Rk��H��Zh����G�M�!��;�z��l��$Ҁ���z�Y���y�я\�)7^{R��A���ҽW��{���X�����������o mM�%����T�
�^��qt��o5V�\#�GNJTcFv�Z�}*�Ӗ�[F��M=���ha��h�y���7bi�k��� ����t>���oB�k���"�����*{U�����v���q5�v�����r����^�u��2�mv��2=P�p![��%��D"{}���z*QŘ�kDI�4v�t�0�9��d	/���k��j�3k�y�����X�_{��w��hhf�`⾙����o,V�r���i��ˆ��M���=�B9�W.U~��mˌ�N����jҞ�B��u�2mw§v��k�"�=<=�-��D��/^5=b�i���� Z���#����}�)'99s� Y��5Y!�H�J�T�G$�{����5;��[sߩ������{LC�g�⟃��6Hi��J��r����h"ݞ	:�h����~���ԘcB���}E!��Y��V�K���G�~�ݾ�������0M�A�t�a�\\��;����t�����2r���W�LPC�c��@�a.��V��b����y�dJb�����4AG�]��|f��۫{�(�O�(n�Bʶ���q��.�P�~4u2�pEu���m��u� ����s0n����<��.���%��P���ʒ_��¾���Ghu;{D
6�2>��𼻹�X��L����;5�d���_�����u?�	�Iz��vXl*&D%eWӶ�2LIj5`���x�Iq����b7�d-m���].�mKl��9�s�<��q(�׼��z̈́5�����t�-ŗ���O[c^�f�����4�!��g���଒�����"aq.�xO�)p�n���n���g,DC>t�}@��sE�ǋͭo��n}T%L�&�52W�Rs��2���}f�!7�Q
�Ê�BO�b�6��x�s���Y@����k�������Ƹ6���d2�R�7*��ڭ̜��U��{?¿-�o��"L�;�(�w��8mo6G9"2F�ܯ<*����/F�N�C�}���5&�� ����o�':�O�
d�l����jOb_AR�ڙI:s�+�	�p�����*���x�-�&�]���A�s��M3y�g����*��>�8�2��I8?'aʬ��^ϴ0`�t��Tl�B��?��� ���K2��Gx8�#�!#����^nA��<\��"%d2�/��\W̆־�����h�=��-{ܲ�Pz�u�_���G�l��S��P���YR!�n�V�lf��l��NU,�c�!�o¬�}�Hxh�|�����Yp3uc��Fu�Z&����`1I2F�2��[�i�KI�{�:���^Ȍ!��KJpޖ�_��(�5X��c˦Ed�$�'�y�g�e��|��V��Y��8z�QX���kF�C����/�8�V��f T�%����җ�55N�j���9�N�w��vX.��E���I��ס@z#�����Z�}缳s���	q�:�:H�jj%�B��,����	"Xp_T�5-r�9������	&A���u�.�
�h0�g��rx;������t�k�WI��
�&��QF§A�����q�|dO�ez�DRsV�
w��ԗ��J���ι�\�"���wi�@%מ�Կ/���G���{�Q7YȪ���[���8*�p5jX���Ǒ���<&��E����C����
	@���1o��솗�wŝ-N��q��5[z(��o5dꞛ9l�2����c���jnz��<9!��}awҚ)B=o�L�E��^��/4i5 �'�P�jݣ.�|�tN�=;XO�gMj�4GPds�M��ޭF�q��\��4~��嫜j�m.
�=��%�9D��3�e'��.��U�蚫<ۉ{f2-��%EL:]�(Vq��p�nV�T���5�!�����eP*�49XDо�F�,�����=�#yYy��>B*��I�d�ް)i�TCǋ<+
e���S���тGƳ�yK�1~�R�޻Մi�a㕎ql�OJ������hac�yn�%3��$#�����[w���-�ͣ���@�C=�)g��˶���V��~�]!��U�٭���:Q�B�����)��=K)d57�=d��h��@�8_�����;����3�P�|rL/�xy����X���&�����2dV�g�*�/���s��Z[�:�h����ugR�ֆU�o'�ԧ@�����!���i���:�]�9�����$;���8K�>T͘���Z���ϒ���/1�O�&�q�X�[Qb���̼E1��la��:��U��ڵz��v˽h
�����;@�ހ��1=���%���a�I\wUO��w�x��[:X=Cy`==���h(,j�v���Σ�[�K��%��S����_.|���:�t�F���a�-�������Y�_T�-U���s��x������l�q�zy>��ق�-:���f�AH��bA����q��ŏZ�&k�Dm���K����p�L)<�7���@����� ��T ���-���� �s���X0T�W���3Y�J[ZyX&s�t�4-�xf #+�q�e�j��x���:q�cDr�4/�Js�0~�+�v³Amp����V��n����"Bį�!i,��XS�A�H�6�{�{7R�F�D��Ȃ⛅k���KM�٤���0@�^,_N*~c���j˫����X�4R�خ�횧�rUp�@��g���(�E��tk&K]F��B*��`�H�-7=��)-׬k	�#��x��
�+�y�������Fd���˨�=����/[إSi���\��������;�$�/��]l�)S��RQM�� 2W���X�r�`�i4(��(o}���<2���yhsU��>b3ˢ�p��b��%.n�lUH�:���YI�zI@4p��
?�֐~��aX��mF��s1P��[&J�G,vQ����~�=�=x�7�A�:7ԑUr��[�칷�%�H�?Ԉ}L��a@�l1�D�F��]��nHʑx;��ߣ��@8��z^ 6߰�8��H�b
(�b�_P��(V�0�
s��eނ��6	D���ka�>��*��H�G�5�7�	}�a�����B��n��V8�W�0�YD��T� ��v(͒�դ�J�P/J?�^wI����A&J)�@8�)�2�p`e�pL��k�ǀ^��rۦ�A��õ�U�~��(�ڽC��%���;!���b���"�k�����z�˙�6b��c+�0�7�^��s�>��U`:����l�C��f�=�<���5���@+��y���/�#0����ণ|�Q���ėq�(�J��rw#-B�Bz�{�ChW�3���.��%��?_9 �}N�sh!����J����w�.�?_���g�7&t'b��`�v�ǥQ�Z������X�������up����%��n�Xg�$�����+]9�u���ܵ�ZCe1��ཪ�/ˈhU�&�y���qᄔ�F7�5#Y�W�1�{��-����D�
�/�G�ZJ�!��v6�B3��z��C?|�a!wXht mߤ{~�I/�{���|x`� �IJ�`q�Q�~B{r�=�MiN=����w}y�T��+B@)ƞ�=%s��Nd�:ˮ����w�!���`���r�i���l<A�����;I�N�Ϛ�����g�O�X�tc+ ozt���<���z[��{�nO�PO���2�!<ĽC�,�B�j2qI��ߔ��y{��Eŕn��P� �L"�Ķ��V@�o��s@h�s��l"cx�V�Y?^e��y�vK��E�Z��� ��F!+/�;t�	*췺C(?�����ۀSO�)S�9�EP7=�����t�: �#���ݿC�W}
���FV��w�A��M��}%�Z� ،&� qD���@>bpvOlvţx��A�N;n�+�0�L��F��}�핃mN���>>o]���L�߹�:�a	6w�-�/(!�ܻ\�es���,#}��sVΓ0�a<�$���Es�]�0vI�S+�|�-��"x7�����R�Z$��K�WCr���������ؓ���u54fF��}��8�=N��t�MC:��K�����iкcw"ӄ�vl�9=V�c�����A�h�!�5���nM9Mx5/�3���k��C�:�Qt�e���G�eK4!P�P�*L�o���%lY��=�߰�W]�ӧ��!�<�hK]T�VcǲP�B�� ��}q��3��U*��� {41"-���Z`�I[�9�/~� �ƎUC8f|�K�	g��L��G��>F�A ��3�@�\\P}i��������C�@Z_�����]�i�� �UE��	V�5�!�
���v�7gR�d��A�Wv��(�~T�/��� ST�r�5$c<:�h��w�B���	�I�pN!o{�X���B��9�ێ�6[�3pgoh`d�|�y�$K��^'jގ@ Ql�������-�$�prҢ��ț�)�C+坜��mc%�vxf����>��ffJ5:�7U�ty�A��S1j_�<\��V��X��:�]o� J�{YR�����U���v�C�F
���?epx���,v;�n�� #�-"H�Q��i���o�*dNRy�]}�?�	��9���H�����)���w(��C��F������c��}>��6v2A3A0��]*�L#:E��Vh<�K���Rrr��J��,Y��{�P,��xBj�GMs���b�ʌ��<+�,w���C���_��h�
�w�tk���=�s-(�6��T�M�:�ZY"Wa��:���Va$��C3#��$��M�:ok۴�/�	ga���Z�6�ǉ� �+}>^��H���4�kĠ̶�W�X�kHX���dgk�Y�Zcل�bg��iJ�Ό�t\{�Z��v��X�e�E�[Vh_��؃'�B�ǮɃ�$.��0ڒ<�n���|�},�L�ѐ���V�{��x�*>��aA���'^�o��T�Xj_��d���� ��G|�Ikb<%/���R�NB�nQ �MJ�}��?O��U�8�V3x�����im'�|Ysȑ� �/M�/}��m�yD��C$����q��j���J,Sa�S3жMn�l������c^�A�<�Yhf����Ƈz�����#@^���Sr AP�`��AU����~/�ƶ����"1X�'�������aDV��P;�E�Z�w�b�>H=@�#���qS7є���+�rg��&Q����f�x�C �w��7՗c��i������G���(Qb]�|O\���u�l�n|�%��� ��E.�Y#�fR¾ϑk�PՐF6�u~u�1x�Ns�mc���r���N��>�i���1��[�L){���� ���n�\nNg�ɽS�\6�f��K�*(�-��;���|ܿG3�]�C`7c��_p8�����Kd�]��ģ�F�l�Vܡ���ݯ#��b/uӥi	��L'� �"�I��͜�i�̏��E��A�J6���3��;��[�w�|�'����`���c���: ��2���M$"){�7!aׄq(�hu-֋�z{���6U�Y9Y�-��4M>�ǽ֠��-�>j 1�BS�F"��SѮ�7M\�u0��:~�/~�*.l��xA�L���:�TDx�+%."y1CF��w9�U���!:�7g:�0ن5����*�C���+��y9A�*�Ҕ�%T�����o���<�1X�ؚ+�[sg� bgx�團���Xt
�u[��R�En���k�W��5��3���72bA�R*�cŰ�(�q�(V0�̐1���:����O{5��wf
��!�}��xC�I��3{�<'Ƽ�HŠ��M�N�%��y�ArJ�)�ą�l{�j�����	7^�i�l}%����;��/��ST?�T쎇2�V���
�9��W5@�A���ZmE6�����c�'��.�I	����a@���=���'��jd=�pԝ|7�A��9��.l��g>5ݣ-����U��:��	I��$;)�L}4����[����'�Nik�����Qb��S�}O!�C� �S�J���)����:d��)��\讷W泽�|�v�3��Z.w��� ����߿`�U��A,��R�������
��Y�&UsO&N
\iAt��~�=j��?a���,с�78!�uyVK_~�I|¥�'�����0�~|���F�zg��*<�U��0��<��҆w�ʅ���\��o�Z��4�R4�Ο�\�3��}���r%�����͂�U��-�����B��Ē�Gh��!��eX|8r�Y8�����ʭg �V�9j���N��6$�rzѹE���~��L���������+9� R���I��"A2�`��x��qU��dz=����i�a�o1���IYB�J��f��Sz.��Y�#u~��`���w��^�X�&k0&FnW_�g�7W�kC��a!_r4����|�e��n��!��LƩ]�%iW5Q����N?��(�S�h��L&��t'�9s7u>�#ht����[i�x[|L/2v�(��/A�H������1�G�r�gk�*yV�B��m�h��kY�L�^��&��ED����!xȯHJ]���w��F�cK`�l�����]�=����W8�DR�o��3O�����&bN�ج؜41�����'8��w�B��ب.�h���y�翔S�#Q9,�𢆘P7�׊�yӈݦ~��Ě �ɋZ���1�Ss�^�ɮm[@J��r�����������R���-�
�ET(h��fN�� 5���٥ް/	m۟;n����msձN�?	�#����rA��gݸ�9�"����?j���lNg���d1K�q�wF�P�RԾ��`�ڕpS䗍����Z��__�h�M��u-�3�*�j�L�)�4J6h��a�;q:iXDX0g;Q���podLDxM��_L��(ά�[�FFU��<)���B'y�|-�+~�O��=�!^�!J|dc��)�f���:Ϫ�g�����!��	�~U�c�� p�pB�M�"�����Lx�4��􍙔�ƨa�,#E�;�����X�M�O�ڒ.��r�}2돱DqXݮ��ځs	����įo2D�+�_��B��oT���
�;�6�f�g�թ�t��4�5%�Ҹ�����Kn����pKi-C�����Y-�T(�%��oU8j��d�շ�\Y����9}_�ۖ�����Pg��<�G�/�|7d�M�IlՂ��������@��?j'_�3R�H�caEYq�oƿ�\oI)Y�1U��V^���+Oj�o�d`�/�(S
g���z�m"��$�A���Bۜ��{��Q�,�_�l:b9?5�'+��7@�[��."�Ѩ?�����,-� E!�cx���!.ho�]�\ݠ�7�&]�Q�P�"���ڱ*K�ae��_kF2]�7h���Ug�*�K?��v:�sSY��� ���QK]]��aU(�*�� RW����<�VH��8�Jp�4sJ������ƍx�x�ݵ��3B{;b�9ʱ��|]=��0$�"3�E� ��4��օ��,}N������4m:�_L���'aA��}�p��q�A�(���#�(�6�EJ�1�5۫GC���勖�+�*�~(W��Do����˵����u�~���q2���׿���^�f�JP�R|�8�-	p��$B�ڃ#TV0[�� ��] = �i/#�
ς��~�Ɩ-Y���������y� �5��uW�k��+���?�]���6&�xDø��\1Ӄ�tkI�'Y��K ȷ�nAX��Qra&�?�������'Q ]�`�J�N�Z�;����g����d �Y	��!�y�YĹ����/`����/Jq޷��NB��	}�^Z��	��16�A`��b�xMK"�ed��,(`��*$�vD�ʹ��y�"ܗ�`���t 9�Y�h>6�M�r��=��)V���7åD��<���/�T�0�q%<�)`Ua�޹8���Y[��j\���G@����e��K��Q��9{������O]��o�`�GL���&l��٣�C>	e@�x{o�ک���[����ӺD �d~��ۤ?����lN���N>ݦȭ(8<ő{vOz1q�i�� 7i�v�3�$ua۱�|��c>��f
g�����z�D��G/ѵ������&4�Ü>�LS��Y��fV0��tQ�?I1\v��[:vD�-Йߙ�Ȕ���vu34]�	0�[� �R��^t��s�
�[�50 ���&+���DOC�L�w�X�|�!�0���#9���(�NH@t���U�h�z'8^E�OU����SMAF�.7����0Vj��//(�#/Q�H�]��)$��M��Aj:��W˄����d�P }
 ����25sk?#�6�"B�\��`��L��Qe睙�xT�o�\��hG(����"߿F��L�oIg�ҷ-2 �QB��*�o_��a�j����j	�țc*2���+��f�F��%[�ƽD�ˑSo|X6�/`+E'�J�x����UUƒJ���ʐm�6�]� ����������;(J�.>��[�@R�� ����D$������_-J���"�����Ւ�*Jy��~��|q�mP=�p�H�S����xܤӿ��o,R���y�e����}vF�Ys�4)�f�����>_�|s@WI+|�s�<�?.)�	i��Ӳe�i(���4չ�?I$ �쓵w�ـw�^:�PC�Dh�x/�^�x���}�1��$&��X�É0�)O��Mc�K�U���<����q@&>���� �;u��O�%��OP %�Ä����/�f��ι��Կ�e+y��D)�g
4�F���f$\�����w{2B����C��޼�ܸ��&R�����>y���_~��2]��m�*�&��]���^�����<b�;��%}�5�=����p���4�:�Ѫ4Bub"�<l=����I'�M�BI�u��J+���JP��Ͼ&3:��V[F��\ͤ�3A�NK���V2���Ss�rn�o���6�S�*�~ۅ4��^s�h$6��(Ձ��{�L2%�m�z�����o�m0�Y�n򇌈�x�+0�K��˝Л틯c�֢����A��=�|[��ı�O��6k��]�|ǟV����
p԰�4���g������wh�f���̍G��I���A��fA)�I�N
x�����̃p�A����s'd^p�0`��y@U����I\�/u��S������b0����d_=��l�ϳ!���V�y����H�]��4i�uV`�j�̋'�!�-@�5����G��3�]V��1�����R�K� �4���|��(N]@�%3w2]�2��x:�?��6��5yA���,��_=��+��������T��Zndf�"	�igO�g��m���8B�N
�af4E�h�޾��i�F-���+�z�Ly��KO;*���Z��$f��dM���c�v�z��tjo�5t�o>�	�C�="��9)8*|��«h�����&��@�Ơ,��PV��}�ˢ ����7r] q�����,������y� ����>��t��)ͱӆ�p��yEe�|�h�e��U��(ȼ�̭s#����؊[�����ǎ��L ���4�j=o-�j1Ǟ�~< �b��]�S����4U͑��]x�g���l��`�|���"�A�k*�0�*hg�̌�����j�����_@E��?X�2�q���3$�&��t��tN`��qK��O�f��D�޹�p�l��m����% O�<n�'#{�:������N�͕oٷ_�t� p�e�;�Q"��J�l���h�G��?#����ʟ�7�B��ޯ��9Ʀ*;���9�����Wڮ6->�X����B!-��`m��U�s_XⰨ�Dj�<�>�	E�%�6�3���&������@Դ;6������pK��'��:�5[ӟ\w�\@�Dr��졩^���V&���q��dؠ��-E�y�CG1�UK��pЖվ��ǜ
��$v)�!�3�Xi�_I�2B�uUΩ���ok�Ӛ���U,��c�����A�&-ǀhg��
�4��-|"�$R�	���pZ�&u�v���L\�`�L.x㷥�IJppLZ�;�뮍@�<
�B�	L�Ŋ�s���m�4t��u|rkV� ��P ��)���o��[�f <Y7��6�U(M\ucB�\����*�.ib�
�k��"_��� ���k�[Y�-٘uF�W���I����a-�6�BR/E>`�@/��	Sy� ���b�)��1�`�%6�rܬ���kY�򷹢x�S(q���1{�#�b��.0���6�@Cߋ���
gǇ	�BW�ݽLR
��"��?�2$lx:(��������`o�U.D(HW��a��k�N��;����H�*D�?;�䏟��B2��r�WS��\���y�r%�ߵ�����y��FP�*�=����5'�Q3��_�?��+W�Ű8�!Bx��@1~9�RNzܼE��ۦ�6��3[ �~�`o9�1{�J�?E�p5���)d�wV��u�\A����C8�Y���&����c��W��4T�!j�<J�����<���j9�i�h6r���cǿQ �C�D9\˒A8��4(gi|�N�XI_�5F��#5*��
_J._�Q�3�l*Ck6?���ݸaÖ&mU*^�Z_�A��ތ�^,�3HT�D��N]�/�>1Ϊ=�]X0�˵NL�� <��SjM�"EѺøsm��o�]��K��po\�:K;)�mg͞hI1e-k�k�8���Ȼ���BKF)��D�eZF�F2l�l� �+��ÿn���'P^��Q#��зܨ�,w��j��1���-�L��x��q���F��?@��:+��֤��OP����/ń��f���=�N�X];�U��W��I�̛;7���q���|ns��I�H? a\.o.W���}3;���!|�@�:֍Rva&lˮ.t,&��A� �rl�DW�=�(r��֥ןV)��ITPLO��Y�j���_�^H���	�m��J��;r|�d<oR�o�aɬ	�+2��Tڟ�(=�b�Ȗ�ݴ��s��Ѻe�����$f@Y�� 
ӆ�k-*���m+�C���jX��~��T����:����>�@>�W����ߪ�B��P�4JMV�~nBit�7�"�����!�8���q�0��R��p(��"(�O�Q�N��c�K)���Gs�wܫҷ��q�;(:�)+fw�m���&�4^h�+9��*���l�z�E3�h(=1%�0�¡�Kzl~�c�2��H��0�(pܟ��Z�(�6����R�g��{���4���u��v����z��G���,v�Q[��:�P�T����ŏ)/A{��q����I�1��K�O���?�ʈ ����o��R��"�,��b	*��E��f&yoK�߅�C��bx|��y��Λ��f8j�* ڬ��bh�|s��҉��4n
�a��,���	�����t�,�����~��j=��W�C�-�����Pd��'�Cţd������J�4��C4��bʋmFЖNo\�Q)�#egc����{SB�0Ǩ�tח���'�ὐ|:A���;6��Ժ�?�Ln��H��*w��j��砃o.������L�tѣI������[I���@$��ᄃ�W�="���F���O����O����4�Lֽ� � sy���:7%*w[x�n]��Q��~DY��Y�/�U���b���<������5��$y��vխl(�*�|W+`�bÁ���y�|����C^hP��W��x�k��`�����(b�ۻ�'-ް�T�����(�@G���Q$1��$�,<�@#�^�� �cc�Z�φ>n�t�[�s�����>��v��AΊ��
���`j�PV�$���NY�V�3"�|+d��&1�*���,{���Bk���(�%��}cҧ)&��ښ��� �53%}�ۊ��+ ��!�r݁8�>���o��o�o����������2�[�;0�s!��U$����X3�W/4V8���Q/�P�F�XE	�H�y6�2
�Wb�x�ޝ�ՠ��ٵ9�[�����Ħ5ځ�����8�r�&`D��s�ϱ�}�ASI��1��d���&�
Kd*ep��K�2�^��h�&Лn�d2���3��X��I�n^�e9%�����P�N����6����:S��t�!�5�Ye����F.f��Q�c���b�$��R�Gx`S�:����v��46T"lI`iI�x1}�.ha���
y� O=S�r�r9iN�b���*Ga$�z���fD�>�lH^�~Rw������vb�V�����,��V��+)*��q��zӞ'��u��D��+?�ʨ*1��O�`��?ͭ5����'��p��,~]�*K)�����������2?�>Dˇ!��Z���C�+��hWTD,tU_�- Ǵ���}�x�ǆ>	xgU��{�Y2���W�����4�|�G
ĩ`�\E���,9|�����'!��(O�?�	�����B��=���\uD"���R)4�mL�#�ji��?w�*᜔�'�XN�djQ5~�l��݋:�D�ĩ�чL?6r��߱�@�� ����\m7�3n�����-�С�J�&���F
��������Q�I�M�J�)�𒡹��f�L��>��Â��A@�0,6�e�iE�$ު�S�ɢקkV1\�D[G�����F'@�epc�X�t��\R�����3_�H>�Z��A`�^�@�fQ����%�{�Ivt4&q;�:�u�L60$M�3Q*���!)xK喩�$�?�c�r�0��_+T[��}����##�{ e�J���7��Ȩ�n?�;<`��<�7�耳�7-�x�Ŕ�$�Ӎ{>�Ηd�Nx����]t���J�*�eHT����A vm�Ӱ"�`y��uu����UR �{P����	�Lt�p���\������Ȉ���)�8v�u�գ���߈�v�o۬��EC��U��E�n4��(F�u��n�)V��D#]��~^d�Z�Fʩ�>�īʡ	2�:�6�`�d�1�V��A�#����r�TX�l��®l��vdd�E)����f��#��r;��Q(�&~N.�e.=�Vl���Ԝ}�F�;vj���Y4����u��n�;�nßpwY��I�PO���Ʒ���s�a �C잌�ڃ�ȩyr�8�P���/ĖKH��iU�}�g�)k[���d�]�6h����2\>\��'�q�a�����H����mO�{�4:��A�U��,7��Ό�//�4I�n<�S7-+��DA8��%�#���Vzm|��A�$oQbfj>Йò�j��ӛU���/GP�K�n�m4���z�V=q�+0B�K9�λMA�Y���bvx^��^0��,���>.��
�T�|EGmr�in�#�@3�n��/xNPi{k�7�":��(*%^�ٟA�i2������[��b���7%7�B��f#LK8���� Q��f���u�W�����V(\=��S��H��� 8����t` 6� �އm���=��-=^�,'��`�
Gf|�@��z,�\�U���VL�ǒ�FU�y�a
*�3b;��M��Z7��q�h��!ӮSg�Nkٵ p7|��HƬ'�o�(�j-���t:�����U��(G)�<�	yT�^&�q�m����8b�Bs���=�L��q�/�������Q���nq̐:\��:�� ��Á��w�E�ވ�Q�_B-��lj�^��-�1�]�zѸ���M�k!������:��r�Df�$A���4�S4;*���}x�1�g�����Šq��������Kw�k	��;�'��a �>�
�ʀ�/�xe���z�s�鎤4}[�c�e~��L�y"~��-���dZ��=!֖)4f�~3���Em3�����Lj�b5��'V�m�<�a����:a��}$D��6a7Zlrj��dةu��S�g}�����n�g%"�9w�qĎU�������YrU��}��*h�k������.�HLvZD��W�X�U�<1�z ����`6�3某^N�ã���J�	���H��MA����8�A�x���ahC��8;�3_�3�mX�q^�
���a����P�Gx�
2��E4�.Z�[�|�Ue�n��3�K[W9US= ��u�����U)��s�Q��Wc�D���c|�,���K�OFI�fQ"hμ�y[���%\L�� ��L(E�V�(�9_�z�
eI�W�I�B3<���W�kA3��
d�wާ,�Ƕ-�x:�Y����/�x ��b��c�¶�1�Z1�5fnFG�]�>����3�I`
��Z���eg�Y��4L��R�8�po�ĩ�S�,��^5s�=��K��i�Pힴ���Y��?;q�HU�K��Ph~�PiX���S	g%�(���`l��m�		��d�vJ���C��@�.&N��J�i{�Y��m�"�#嬈c�bKh��b���Q#w��1���F���֪~kL��Q��!ݣ&�Y�z��
)�RQ�ʹ�8GY�[1O3�$��Pj(wdП�L�������AH�Reї�*�[,;W��r���)�������)f��-ݶϽ>(�S(���h{�0T�5��|�B�y=z�ܱ�<N�߃�<R�����h��T�	�t�N�t1o[i�z6U���jI�1@��&��ζh|^���A��Arњ�aG����UD y}���tq�"z�3�P�����9m{b�.q�0P�,)���'��E��#
Q#�#��.�9|���
k�J����
�[	�~9Ļ����|+�S�w�|�,g[�Z��`�����K�b=�O�94��C��ʈ�W�4�1`��;����������pG�C,�yhai�';ص~o7i�S�+#�ժ�$�,xрB�����ѱ'��{�E�0���6yb�l�R���Ve6����Ddk� ��EH2F%�G�1^�_���I���}�D�zmNf�{����n�F�}0%�s�&�g��#f��!!U��؊�<=�:"TY�e�Km�ɉc��a�$�{W'���Yj��Ϯ�L��,���H�qG�:��j��|���[�����ui�ě��%3f�^+\�)�z�8q'�H����y�o����Q+�!�}��ԅR����m���\���<��A!����׎�.�V��~] B�l��mU����]�U�ڃ�������	G�Q>���a���ٻ�������Q�6�H.�ł�O���R��^�/ҥMD�13��5ͼ,%�92�o(�WI��Ʒb���]g�s;{�3�J ��t|�=?�9�(�Y@��o���oeV�x����\_[�c����A\ ��:���#��|�Tl�f��e�ˎ0	}�=B���:)�-f�"��qd�]�w{��Q��θ_�m03�����pKІ��pF��;�>��d�5̦�,,���y�*CI\��a��〼ݩ�[�hd��f(��#@H���g�0�.�[��Μ�]S��7�k$�$���a�u'�xV}���:e�7�	�׮B�����I3������������X�Y����"��~�qV�2�"�fx��PyU� Mhx� J}]����$�
J�S�cL����١��!B��jo~��oN�&F�p]P����|ZX\�O5CE1��g��'���J�E���[����4�������s��(�>��ճ�}t{�w���}2{I:¡������M&�U�n�eF�n�ZaFi9�'��ڌ��!m8��u��?	���{i'���P�e�;?�����C���rɨ��̍��1�b,���o��������@��\�U]�O!V8��7���E�'�:hi�t����_��x^��G   �KWG�����Zf1�o�Dq6��NЮ� >��qA��ʨ]6��fEj�����j,����3�H�ޡ�����OS��8��4�d���!L���p�;Z��{7�ɻ�,�������.��9�In������a�ȟ��`O��:�|�Oȅă��1��<��`3�`�Ms�^���b7����ۄ��*�E��2�u��v{L�b�,��$4R�<*����q��P*���!<�Ζ�p!?7/�J�N=>�A��&%?ծ��[7���D^H,��cWgA*�ޮ�l�W�Џ�x�U
��V�f.�!��
�x5ť,��WR��[�Wn�dS�W�����bfw�&q�aZ�C����|ù��q�bM� v8�{ĉ�N-p���uƤ��3�'�`�?(��	ߨ�C����"38ӒH�z�ͯ�|����ܹ�U戚� ߩ�ua��e�hM��]���D���)��XGsp�)T*	�Wj�N&k�nen�c�Y&�b����8&�BFf���Ԭ9���l�l�(��x,ȳ��,�.��#�x���#;�qK�<G��������NXh��ՉE[|^B��M��$��o�����B�ٽ&�0#����7��P��6�_g�y��>�R�)рә6^U�2�N��=U"��N ���+N��!��Ÿ
Z;T� �tpl�-�lg�ɾ\�N�6��B7tX}.�D	t��i�S`}uJ˾�����Yk
 �s��ܮ�N=�9rR��5e�AP��x��@����Q�������#"�\��3�t��ǐ��LAX(��ނ~W�l�-��9���p�T�z�w�(�pP���Rf����U݌�rY��t��p���F��R�\[*4A����dq��P�6x��=,'Ɗ)�3��E���R#K��m�vEo���I�RW��m��ZN���y����`�h_���~p�d5l|���C�H�=�oVH���E4���T���tf���H�����	�[E�������׫�����n@	["�-�;�1Nɭ�Y���KŹZ�(�_���Z���*k��α������,_�U�X��!$�{���Û��nӊ��t��-s4>O#�� �	�0+�6��ʴ(WZs���E�11lVWu�R�ؙ�n��U��&~wƺ0��M�����.��$b�����0�ER������]k�1�3 ������]����I�劏z�'%�.�/�@W�(�OKT����9p׻rD�"�j�ܗu���a��$5t�@�CِP�S�;�&�o�f·�@rr;g���K���%���D��Г3;�T�?���f�ës�T����A��4x&�_Z����y��X	���Y�zՀ�Z�������pz,P��p& o3��zA��),+Y��S�(y�(l5�@ݏ�7w!s�\]�XKp�q��W;��w
����{ܳ�Hu��n�wy7����O�l{�/�,ޯ�A����r_:���۠y��C��n&s,�]NvU����{���9��~'�3�H��$g����d�;�=����U|��l�j`-������������Ho0���Hzly@=T�λ{[��<���<7(0Lȱ��%]%j����7"��>������v1f7��0��
T~(ܥ�t������Q���c���hg�R+^`��d�J�8�k�?��4�ί�k�<a�od�'~��12[����'�/#G�lO�G�s��低	+�,V��2.�=$��E��_9�RԆ�[-�R�BS�yて	(�����HKA+̧���=�n����S�T	_0��YQ)N��W.MY��{�$���m��i1��z��mI�Ǟ��S�Ú����-�!9y*j��
�9�2De��>�����WS�r�x=�\@�Ƕ�1� {,M����m^��*��z�m	������������[k�I���"��.��Lpk?i���c�r�I�yD��X�V�����������d��l$W���Y$�v��A���!\�d-I,����T	�h^��v�v����"�<��F2iD�8+��e��V��t	���)�b��`%�|����(�ǿ��y�+��h�ZV��Z���8�X��3�\��ӗ08����P3ї��<on�����"�}\��ۤ(i�X��@/�ml!V$���3�1�X��n���/�.+k�ړU�QS
+̓u*O]Ԃ,�ئC3���ғpy]@64\�4����&�,BR�]&��!�[=�����������]Z���nA������h�����0�t���H�6V�@�^��QuJRb���k��>Q��H�\!�{f���PǼE�E5z�5J*����¾Vfm�Eq9�V�GmL��a0,�p$[5`�%G��E][�������<-s���kqϫx8Z�A9Ig�)���z��W��K���e��(u�2�#h���F>��FW��V�sM�`5�R��I��8I�c�ԌժB�7�U���V1��`|턲C�W|R�$�؞�+�tIs4����qW��=mO�����عzP��w���E��e���O��V�\������o�u��d�_�~������j��b���&�L�$�n����c	�Bƣԟ �rr��[t�?�Z�>n+n���D�Y�k��.@����b����PV}�'��)����~\8ǻ�1�Ju��!��g�<�m�jy�����K�,&y*qf��k	&o�pge�  �/J�u2�X�Eu�>�B�q���k�xI��x�������ٺ�َ�z� F<9��=�G���W�<\�huq�5���F(T�>�1mf[i��0�q8_#�1��Չ�H����������AK���Z���v�~�1d�k�.������Hl⑊�x�\N
���f�� �}J/θEL���g���0S��Y�X�(晊s�"����B��BB/)f�}��#�KڣG��¯Lu�mA{М��nhe��
��OC8����16�2�e3��y��p�e����%�¶R+JE�Ӽ�F o�7!��§�]��Dл�����P1����?�6��J;2��g���u�$�~Q�@�ѥ
��v�Sb��TΊ��O;�L�a?�e��*�(<�6�~"���#-EU��8��(0�"�4�ءXy+�N��U�TS@E� �[6!����yb�U����X����3��9��>^f�}"�G��3��Jď(ˍS���5f����E��K��]�ե�_(ڨ�_PS�Y-kG+���sD����t)��F+*(�V��Z�٥E�E�r��6 U�0���WP��
�x�ψj�Z�5eڎAfk�g����hк����?J,�{�cö�5�:l�ze���؎:x��Sk�*9��)G}��vABU��L)���;��D�i*�Q_r��C�\v;��ǆ�?�˔�'�\`�N4.bv��N�s}K�;��B��� ��]k/��O��d�*Ê�����`�V�	Ƒd�*����e�2S�s�S"�t�X�+��R�}|�7~5*��+/Ե�����ښ��W�9����s���|��( �W�������O��)PD�x;4��
�~Z�sr�d�9Z h��=ԛ"UW*y�]�'��
E�W��<���5$[#Ȋ�\]sf[7�S���||?Ұ�k/=~g`�c�A	ݬ�FN��U,��k����)y3T��5r����T�s%���8�H4����Z�d������e��O)�+�>dL���#y�I��Y���(�|��U��O�Ѳ� �S��� "/j��(�u�~��({bK+��9�~�N�޶ 	�.��E��7�F�y+�S��'�e,ټ�]�	�q���|F\d/:3����q,İ�L�ո��/����^��q�1�kOr����aj�)�p��"уѧY�[�w_�lM0>���3X�B:������+j��Vr�2[/x�"��~"CLs������mf�&.xUq���A�[�&�0��}�]��'�;��尖�##��^��� ���ѣ��M2iٖ.��>���k����3�\:<W�LA����J���$�b��h�OԢ|��	D�J5v&�PM�D�����'s?��u�ȫ��>a�j��h��V)+7Z��.;]�%��7�$��Y���|�qޙCi�Ta��ιQ9�P�4 �{�)b;8��� ��x��?@2`Ӈ�����CR��@:�����VA�kZ��Ào%�������Ԍ/� u���V6�ʫ,-��&�`����ܾ�.�5|tE�,l��x��7��ݺU���'� �r��[Ny��1���g"���!:L���C�1x�	�N�\��Ǥk���������śyr�N�q�9� g��e"�-\Iy�f�D�>m��9��[�g�_�?��0e̤��n�FӦ���].+�0ml�9؝�Hh��])	��,������)\�<>����_F�g��+ � �SOd�M	���hP����,W� i�-I 荷\����`ݻ\���G�g64�wql��X�n��Fk^��`j*Ul��O§-���\��lCx;<��ef,�;i-l+�}Pi�?Px�}��?���0�d:�9�/ @S��=��[�7oM���X�̣1����O(��JC9�����b�����n��a?�c� qJj�"���f�g#��q�S��	�(�hƩ���\����>"Ӻ��6N�����������G�OƓ�33��1�p�M�|��R9R��#}4n��p�KH����d>�)��*k�c���c�^�UF��P��e�۵EW)�f���~�Q�6�
��|NC\g{n�Tޛ��o��]�^:�;`֩/���i��q�Uӊ3@�@A?�����#B�����&3���6hH<c���r�,�Q"1��IKv:�Ǉy��[��a�%��i�fZ=7��BV̳���FpQm��J��Zw�d�NcQ�9�4�'e�aN"��ٳ�їR �K���7` -�Ī�^ѮI��ۡ�tr9�D�@��ƺ���Wt��ȅYD_��[��w��Դ�w���O	6D�+us���7�}c\𼠾d��Р����ގ5��́��F�l�%�*�vʋ�9a����I����W������[�by��!���GX��8�?���Pu�@X�a�<jiHE�S*��}��1K��y�[����I�	H��9�7���.�C?ė��4�
�IҺ����x5$��h��g���5*��O��N�����̀���f���]���+���qi1�7�Rw��h��
+Ɂ���ѱ�(@͗84tcXL�$�o�,�Kw
��$D���cGj����W7�O]����a��^0ѐ�Dov����T�ә�,�9h�AT.��΍�&���ig��oO�o���򕰪��v'��`�������c��Fr}M�"��\4�mMCN��r�K��D�m�{7oQ��N�|ᜧ),��D�&2����)U��DSF\i g��D[��}V�#䦃��@�՗� F��g�n�9����>���3o�uuQ�E@'k�f�nB>%��s*��>�Pхi>*[~��qmQ2f���H��V:�!j�AU�ٚ��
�&L����:1]�7iA�Z;S{/��?���*���z�C�ǳc�ER��Ff���#�}�l�4?�Hݼ��o�Ez�`j����d&��)����):3>�C�?��h�a=m �Esi�~k����8Z���NP�u%�Y��,�$�OX��`v����$U��X=�3O�R���+nʮ>�FZ'��;�4�P�W�JL��;��њ"M�JB���̞x��@pN���n����v���`�szOF�&gyQ�1�>ȋ��w'��N��$p�f�P�G�c6��2Rg����O/T*�� �c�>ޛ%:�m�S����X�hXZ6�$ z�fs(YH���VoN->�_����3Ő�C_�VS:"p�ς�����R0�p(4���}$��D����/��]��D�#8y{a�\Vش�a�Q��y�ୄ��ԛݩH�P�@�����_އ�� ��+T�%�r&��G|/(��e֢����yN��I.d2�����0����ڲmHNPRoI'D�s�̩����� W!�*C�Gm���ٱ��U����<�fj�:�t�F��x�,�{j�H�1y�����3�^��DX���NIFQϰ�ɹw�2U>ǻ-�C����E��ā�{<�����jR⑃���a��"�υ1A�(+��q�oa�Wvqީ&\�-V���U��6Z�R���-�\�p���7k�	dx:Ώ	�=�����7p=�v��ܜ����o�!e6���66E+�h X8oF.�CL�z-�RJ��>�HGZ��W���n�8S�����LSc��s���6�(�~?�	�
�+�vd���|-t&SE��M�(�/״����m��$Fiw�T�%�#����w�������<ݛڠEc����1"�e�n2�CSޝ�*N*�
�=j�x0������ӊ.X�D���E�Dʢ�����FB��7�z�o�ʋ�qZVE�b_4	ilc� t�#%��K=�7�R�w:�$����G��{ܦ����D3(�,t=�q��n�α��b"!�HST�x%�X��.K��r�C_)_�>^�gA��W��]��Aۡ����΀�7���R���U���Ȍ�\#Al��Y�Pimo��e|��2�y�6�:�ġ�)�RJ-8�~��)�+�K����*9`�j�#��H��s���۔��H4���1�H؎��7�S�ǈ!������ʫ�T�J���*��r;��c���.eA�&�Н6}P��0`���y3�t�_7��)vsc�'�9����B�'RYA�l1bOv�X�ـ&y�R��a"[^4j�s�l`�K�!�&m|���}C��6�Jp"Ej��{|hRp]�t��ңA������SV��N1]���2��������c�I:]Ψ�r(i4�S*z("�����w��n��Au�d�sC
�n%_o��p
�����̝�:	yq�]8�!Rdn��0�-Q�H"������KSu`I*2�	(��;���>������|�8�ߣ�I�2��Z��	�F�yN'>\�Չ,g`���ބHW�b�fX���8٣3Ť�V���o0
T��t�O&pM�D

~̿���Q��¯7��^�#_[��f���-��jt��Q�9}|��ı�s-�$n�����xQ�{��9�Wx�'�\�O�^�O� � ����p؀�.;O�-h�t�Oc�V*��K~>~�d���$X
�k���H����3��&
y�P�3ՠ����V�L*A���5��Z���$�9Ob�-ѡ���Oߍ�RȢx��6SE�4 ��KH!����̘G#@�eV9�|�l������N3�LN)�t;�ifj 8������"9\2pNQ� ����@݂�]Z�iO`x"��
f�T�K�߻��|@1������(�cU�퐑YI�bʠ�nn�I=������H��s�A=煊X��%�F�9H�]����Q%��B���L۔�����;
�-Li�"�%Wd���\��!U �^�Ŕ�#�%�[��>�mI��C����9�d�c��7�4���h�K�z����������X��k�ʷT�MN���וk5XЗ Լq؛��N�����\� c�{{�oj�R��#	y;�_�4գ��#vE8WuSb��D��l��AC�&�F0U�Q˂j�/b}�y�j�۶�] ��"m藪������v
�vwf��a��;)�>��!�"_�-�@�S�
U�K㢆;$�E�PI���I0��� ��nX�*��|��l��e�ƥ�ե��}� �I�N
k�x���:�뭛�Ց��/>���L_�b����k'�:�oAX���o�y���
�	���+����֭�<��� V��;���s�7�A��ߎ�$H�а3.�zc~�3�/���В��MK Oee���Ϛ O߀�}"�B�s�qԶ7�
'FN/9XO�V[gd��:�b�a+@J����t.�T�B��5r���~-J���3�x@�v�S�0������X��R2���y�WNOI�RG�B.r�A�2<I� D#���x�,H����í8��u//Pr�r��M.S��d��׾��!1�%��|��8g���w`	V��W�7O�;
dޛ�Y�{w'�}RC�ob6ꑒ����5��;�5�iY2��A���������Z��&�-��C�y�o�5����F��Ő~�H��?:/I�*�)��"&o��a]��)�Թ�+�(KK�T����q*�$���>_�B��*��^���&O�և,Y�{p[�T��ɝΤV'z�iо�1���i���pty�s���qE�t�b�O"s~��"��R�b0 ́�>�Q��U����LpԎD�=#8�p����yL����q�+��sD<v��daV�:�j-Lf�Z�E�Y����WV��d��4N�#'��It7v@M�`�ӧ6|ؾ:�ڷ��R/`7�=I"�����Ǚ���G�`1�0�[�/��q�A��@��A�w�UO,_�^*;l�$���u�������؇�p�5-[��͒4�Hy|�I��[�*m����;��"��`Ԑq�z�_pS-rlY|�(7�q!�;{`Q���^�@I�OV��yuMl�! wJS����q�ez�͙1�w��!��^�b�!_,
�Tb=";���R�Q@�s$p�T�N�
_tQ�� Z��VV�p�&�D��d)�gaS�������2�(#F�iT阍^����|{�X����B�3O
��e�aenGM�PJC��x���e+CHu�F@��E��b��#q�Q�:*��j��	�j,���m�{De�M�뭱�[�W+�� ��t$���zc4܀��h��W�!GvV�)�Bv%�M��2�M���P�2n�3,uTE尾av��ʅ�h��2Jz��Z����_<��}ҳ1��R�]D���G��z΍ ���.�*w1s7�<�]�s�d0"���\`�/��2�C�q㰝�S�=�"h+����d.K���9]��,Hx��EBq�S&qmn꽯��=��n�FJ���G�W�K#�{y@^�߸*�t_�{�ރb �~��i�"0f��Bj��LFiMJB���T8y�\]��드���Q�i�JF�r�O.�/��i!/N�:��N����Z����_�`���9f�7�aɡ}�AA��	�|��V �خ8C�ڮZ���H��ߟ����%Sy;�ݢ�}Z(�P����v��B^��,�m�H�������|o{��1����%�J5'x���@r99�y_+9a{�����1�!M���w��p�P��?��'"�)`�Go���[��*�9��3g1_���k�e�3.�F�nV�g�6��sk��Ou^���N�pA�%�����E��*m����]��~A���0>����1��9}���>�����J]�@N�d��/;������.w�A@K�:% m��
�$2EO¶�!�����r�N(��J��w�`TL���-t(�=.ao�87.,6��&}Z�?����b	-g�%~��J�ܴ�DT%��N~����({:~�1V�MaLp��ِ�"�3�|�7xy�mU��r�v6��_1qk>&=W��L�ZNT=pa$njI ���Rg1i�J�(��S�P�W����S{�cˤ����nXgM�`���Xl@�a_tY�V�c�T��Ֆݧ�B�u��]��X7#yjșH����/M�� 1��Ǣ�*A!�0�J㠑��*�lbN����2}Z�t��U����?�wg!�"4!{S�C�i����hO�#K�ְy���[w�=�g�܌&����k��$�Q������|���z��2-�Tm�����(_Dv��%I�	4M�7#�,(���>��V�ӽ�F�@�i����i��-�A��腵��`Ȣ	�W�'�9�QιT.h�6:�>���ٝa�\�K".��A�dX���G�m<��_���v�"�AKO���-DY#�|}��^����WO�	ː��$�Ծ25*Ɉ������N���W(�+����Z= O���|=w%N���d	XN�^�p	KDgzY��z�!�VGv��{�fcn0���j)զ������e�F���[�b
���y\1l�<yB�+�������o��N�o�ܑ����=�?����}H�Z�r6G;CYlm���q!��^�WEb�0�[o�y
k
�,U��c��p̋��P��-��夥s$��9#�xw��^��p�����?�d��>5��`���b�\{�<��qA#�c%,�f=q������9SyH��<*�9�BCڷ,���^u(�؎���OK'J_?ΧnQ㾴D�r��K�h�����M�>ud3�
	��*�*�طcT�uz��M`k���q��h��&��ޤ��L��#����� At���+�l�8�^=�k#'���畣d�b �U�?j���+�nN�P�{{�G�C��Aí��hnƀ�oH������.�J��ٴ�&e>v��[�6�2�ژRI�2Շ��x�Ps�D�}�y��	ԭ9�^]�כ�m�-C*��C�<��6��T�b�󙼍�n�11`{�T%���Õ�N����*��]������Eo��+���撙�
+��zf,To��,y�W����y��C̹��3i#�9���(�S�+���Z�$V����Y?��ޯ�C�V"�K�=�
�]�d�!�����mq�K����Hm��	����B�>�خ�5��ʻC���6w=�!t��A�SwW$�^y��D� ��U���A����L����V�`�ɐ/,���@0?�y����Q�Q*�ȗ7��,�g7�(���=9M��r����2��&	�7��	0����!)x����i�U����)�YjZFf$w���(���p��vHO�����0�+��<Uh�i��+@Kȉ#V��O�a*��ֲ���z��S���rF^F���<s��'f���tGkwԌ �n��ʹЌW�t.�($`�#q��eo�J��Kf e=�1���������IC¸4K�y]��	LY��ڶ�P!��^H��6�F�t��
c��W'�u���Y�TpO����U�yp_�m0��ux:6}%�98M�q���})%��yA3��w_K��vT�,;c�j1�Ҏ�]���V�)���Ɛ=�����R���	�hx1(?�B�V��N���.�����wb2-��y��g���ǀ�v��<3Y%�QLv<���w�>��M�O���r8x���&Q,��?�^��Jm;	/{��=F)��i��_�ǽ���](eym�'��,IBCFz�gc8�/4���i�Kqf�@��;�g�ۮ�(��2VB7[�7������4��m�y���"�3����ַ۲H#�FhLS(�u����Ȑ�9�>Ӷ�K
'`m�P�K �CuoY�U��8x�X�y	���Цg�܇E궁�7(p�����o�w�&7 ��8�!�P��"N����mH���q����%==E����&-�<Z�=�E��Oz:F7Ȁ��u�@��f�0��fj��.��:,�����N�Q�.�T��y!zG׭�'솊T�X��#K�$'���� � 0�YvRæM9ь�i'��]��&y����X���/5I���A2 :�j�oM�7?G�<�/���T��D�-�׺�bU����A����Mq֖���z�4������O�J��O����ڀ\MJ3�vьV"iQ������i�Ed�=jl%&��^^��!G(��;a�a��
�m7j#�Pl5m�Հ�Z(T����WL3�l��)�����s���*EUӁ1�qlhԤ�)��qڹ!@f�	!�8�e�ʼO�6Lv��lY���k��B�$H��C�f��|�z�w�E�\�s���Ud ��]���w^�]�=�a���=ٚ
�*�ȫ�(���IhP�Y�[5/�Vէ�A�N6E_�b������`k(|e�+,|�O��X��ڊ�Z���ɜ��ߐ��O�΅��	���Wxk�����z�֎f#L�,-r4U/���LM_�Z|���
�P�#*G�8�Q5Wl�s0ϋ=��a�@/s�XNӰS4�օ���W�3<�X6���Ͳw�;zʢ�7���U�ha_��k�4���1�${ �y���{���N��e\m����X�l�c:��p�)��eVƭ�����l{C��&��ZA�5�v�u�cXRx�F#
��cQ16a!ڴo�?�~��	.�vfgC�����:)�qC���±e���q�o_�iV�*8Pt�.]�C@
�T΁°S�b38�p�)����7���9�-9�	�����ZM�qQ��
����ڮ
�r���9��hV�G�;�t�˿  �b�%j ���<[��,dRD�+۔��g�����>�G� �YPy;��j�>v��k����ϥ>���p|�t�N��+D�R��0�u�<0}R�� +v���p����a�8��xc�l����KTB���>�?���f�mI���^E����O��D������7Y�@�͆��w�q��5���(2ӧ��p�|���8i�I���l����_9�}ki���!j��yk�F)ߨfI�
�ƻ���,����'��w���Y��`wAx״x�n�R��0D��SBc�*�7gΓ� o��x�ߋ�q�G����������N���g>O��{c`�%�R�ۗzy�ύez!�M$��w���4�5wb�߃��v]���b���*Q�TS\��b��S.G���m�\'�.m`D�0����wl$�GM�E�Z{�t�0�����D>	�#��o s��1s�C����N���?��Mi^�����^�]�y��lv���	��r���s�����4�Hy"7��Y#]�ƪ��z�-賲]G�F2��csm��W��{�'�od�b�����p~Ʒ����/����Q��aX����el5>�9_��u,:oH'T�+T���������S&���]4�����_��U�w��Ǻ�shM�U^a]W�������Pz��-�m��}���V�P��d�^_���1Ԟ��n��G��`O�sCV�v���y���Ȟ�Cs��QgY�y��j�u�pl�'�<���mެbJ���h�̊�^g��]�:]�66� ��4j�+ ����K.GB�Ǻ���H����fRH�>* K?M
����K��s��@�$�@���������*��	�>
�e!��M*.O����2��Jh����iS%�#?4z�kN��3����O,��*�~�9�I����g簠Y���Ǵ�i.3��4;���ܚ��>���͚��i7��j��nB��y�Ĕ��߫�q�69_��(`3���'�ﺘU0%��[C,ߏ��cp~���Ws�y˗*^;�"��ҍ7zɡ�!�bT83��U�N���o�63�$����݇������|0�ٴ������M�>��9�R��n$���%��u��_�����N�X�E~���6�:��"�k+�����{�#����/��~����~�� ȵ��I��,>A�k�J��-lZ1�aJM3|jI��^��9��4��d,����g�(�<=Bolua�<��W�L�Q�{_�1*2-,������y�Pސ&cgl�֘�^xM=��L���.щ��/{�^��o��}c��oK*�~(zSL�V�#pM��6A����> �'`�~��+�2Kɜ@�@ۤ��; �vrr�|��{բl+4
Z���ɒ������l�)}� `���\6�|3]����$Y��?�|��7�SV+����.��G�4����&��TqFwCf�9/F#������j)��P-w����׉�OTR�S�a���!�!���U�O���M�w.��y��9��G@�@1���y�ׁ@Fx��Sq��HAO�Y�U̪�@�,�Џ��.W)���y���r3)��!L0g�|����{=z� ������!1FZh�X��A�pTWZ���R>?́��Cx��P<��5��Db��o�m+(L��d�Ƈ�,���Ǹ=����z4s� ���N謓��#�O���-z�\��@�0|�^����.�8&K,OÉ!6�'<b�UY2�Z#~�Eshb��LY�g��<?�����K��"MpOv1S�hj�������
��-�,cW�~9���zy�@��Y�qH\�hL�t�U�YgϾ|-�&PhwG����k��#1�WN�@�cY�ƣڿ!�������	��a��������Bk�zio�+�̽;CK%lqb��Q���a�4��q�B�ol�]��ރ�z�m��ABCe��qn�JI?���O�o��4��g���:�:��)�YUNZ�1� qv�?����C���#ڧ����G�U��ٗd,��U	��'/+C�Э[I�e�.( .���T⤴>��7�Y��{�g���I��|���q�	Yy*B��p��k;��['I}c�dDir2>$��09(�?bkP=�L{oh�;w�X�d�
U0.!5Tɫ��F�)�}��S��@"�-�6]��ޡ���]�y���^)?�Ӓ�&��"iN�R�-R�Ԥɡ�[�k`[>��3ȭ{-i�,d�����N��$XN#�1��;J9� B$a�{���ź�	��tL6t[���7k)d��)����<O��I�c6&��;Ό����Ir,U�JB�.�O~5�vm
"�x�Ѡ����^*4<�q����&IVW�����/�SS���	��!�p�Y�#��] �vc�"E���&M9�����@�
���E��S�~ӯb�ܲ���`]1)��k9W�����+Ћ�L��P�B�Q/m����^h���f� �d=��Ac�����y鏒�t�a�LѰ؃����RnC����y�E� p/��pjmB�,�#-C��v�>1���Б3�E����A���
��}��_K4�a{Z�je�t;`7�O�QC�A4`?���U|��Q͖V`�D�.�X(�v�ݱ������,�`C"P�Z�T��!��+v	���'�^[�%�Gf����)Nwn��M�h�ޯ��F�IP��?�{�F���y�`T}�6���5��vHy�g|_';���p;�<�9���e=��؆�S���Y�/��MB�sP��In��N}���P{��XE_�ޞ�������E���;�o0?m������j���9�E��-� 8�m�o����39j0�N��$�оJL�b�͕H>�!<�^��������bR� \�]��"�6B�1���V���u���/�[��~���=�#������H�����rB�����WR���t\�$^�A�Y,�a��:��L��t��)�!���N ����og�v|���b(?�=?��~CȾ����7q,U�S��A�N��ZϏ6���}�!?t�zlU�ܼ-�N���AA:��q�?�.|O�[bF�}f�I�Ї����G�hN�o�U%(7�a	��fOs?z�?a��R�!��@����B�C@/�����w�r����z^��a�)U��>���|�]5 kw����K�r��R�y-9~����d)1a��(P4?%��Q�A1����5�χ������&�/X@p�^��}�Hn=[D�r�R�.yɲ2���Ĉ�:hy~��g?ꈱ6�H�6J7��^b�7�/,��a92���|�>�s��F��AA8d�<�V�sI��`�?�M���)��0���ii�s/���R-�q��L,�������f,��
���I�ݾ��	�v#L���bxS��_�O��tplvw���g��zܘWQV�OQ+�@+�Gg�F���g��O* l=	yW�̻:t-Ï�;MO�P")���-n��j���Ë�����=��Y�R��ވ�5��9��9z�BȱxigOgl����������C�U`�B%�EU�j�h�	J��X������`Mg�����r���W��Sc�v��u���!&�S��"�vp�^y�64�1����P����{Z�uNf�N�b������*x�Bfu���U(&�g�c~�T�K���D�H1�
�8>l��|<<����хܹ)&a�9�=�'��z�R���{r$���g��6�,vQ�-'���7v��غܼ�t_�0��6��vMs7hş���J:,��;UW��:�-Tp=SRz{�����)�u�I��������LB�(k���D|�Y�=�a�tg��g���?�tóY�gޘ$�dq��/
?}h�R6�,>�4���ǌ�q,�*6ǁ�A��K�$m�Ċ��%�<�,N㓡`ƫx��Ub���4 c�Q��_2���]A)s+\]3��ۛxkT޾��B'�K�N=�!C�S��A�Y��յ���h0x�t�+]�.�犎�5�mZU?m��<f�7�+�0���.y3ћ��t�/���g�JGq�s��[hR)�A��E 0!y�/'l'^a���^dz��Ԩ�A�MBڗ�3c(t}]�.��1˷���V[Eo����E����?�NQ�~��o���ّ�"��\q`e�Ӽ6������� 2�lD�E�i�	��C�@[�|Kxo[��d��N���Yҍᖮ�c$9l����޲,X"P8:�/���*�u�@p��rL����Uj{�����C�J{X�a��	^��Jj��˗�o�j�c3���)Z
��knr��L���m���m	�:�U碻���M3#$w5�M�zE>�5����T�bm�<�Ib��Yf$|S.7��A
�;1�4}��	[H�c�a�|`�X�v��]M���p2�u��R����0�\�76���{�Ǫ�}hMh"����D�N�anG�Vk�@C����0�'������>��M4�seL�d�������^
���E>��+�
�h��K��+��a]�/���W�����rj�0<�� G՛��(��G�E&�-n��������ܖ����"k�T���s���O֠�K��3p��h���7ӂ�nc����BV��z�
�ŠN�T�Ǧ6��t�mb��^x�d�I�`�J�\.�����dX��a��DM�Qc5�S���V>hU� י��K �nt�&?�����bĨ�C��T���*�MuX��f��,=�%8���1E�����T��&�08�<\��Yb�]g���x��[��t��Y~��]`TL�R�VHeM��u'���M>6m��oC ^<�$�����5࢓D�r�����jf
��q]��uh{_3+dax?��f&(�,T+
���\3cx{��R����*a{�e��C�a�V|\DU�iZ�n���>%�z[m�r@�"�+R*2�ݞ�r���\J�ZX��F�A"����OuC�;,FgH�%9%Zx 6Uub�2�z&D���� `X�}6�4vo���~�i�eFjŉ�CH��̔Ǭ�c<��3b���Q��Hi��_�y6��i�ܾ�'��S��ˈk�)33��va*J��$\�W���J�8�9Y�J��·j�{��u�f��^d��7��,1(^�Vx��i��������:�={���0��,P_,���,�-d�>S�4���L�5G�}�h�|6�؅���X*�~��x*m>H.��iM�	A�V�je��'�]�T�v-��[�c%1㩯�<�nT��	�����MNvA��ʊ����1��:�!?6d6�q��Y��R�{�^�oʑ{� ���ٚ���t�����хnĤ/�D=�l��~#�@���7a*t
Ob�m��Ǟ�q��ӂ�������;P3f�e�K>��=�^Z����_='��X�դ�`h5�>͹;�Jye:q�8�1/�O�w�����o`��|({q"���m׌�+!r�����Y��[��g�k��Ї�B}?���LQ{�����;p&�I��K��Z;�P@�Ф��Y+�O`�"c�o�R���z�$r2�.�B����7˴g��Ѻ�;l�e��wB~�!�ّ0�kk9�r������$P���;�]g"*����]��� W�,��YJ�p��
Kڐ�`�MB��\u����.�zk���ޅ_lɈ���ӧ]MV�`�4U����;/;�>����E�����c%�>c�nU�ŌO܃�y��H�U�����J��Bљ���ืRg:;�AP�0teK��x��1�E����56�oUYGM�BP��k���t.�N���;�8z+x/��[@