��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� rā�SZ )����C.��&0C]�-��[�3�-���+��պݣ�k�J�vo`�A�����f����u�X���v�=�а���]Q�Wۿ�߸�=_Q�X����j>��Zw�K��SvX��ƥ.���#�����Z�0���#7{��\S$��@1I�QX~TQ�E��db����۰� ���>0�%�9�j汈��}��1� ��2���h�G��SeY�a���	'<x�p��k�H`�H�j^y�0�s�78+���ֳ�`�R3dW��_��{p[�?$�s0��#�zS�_��bH
�c�p�IL7]� |����Q�� ��Rr���=��E즕2%�����`�^��l�q-�]�p��jf��Ӽ-f%H���ȳ�>��+���M�71��4_�) 3�46h�rb�J�W� k�h~K0�>P$�_n)���5�r�j��W�J&޴o��$>��6��ŀ�;A~<6P��K�~��f��*I
�Z��}`q���ApC��n���g���3��-�іrO�mF���,�$��@�BI�q�}��Ȥ֐����î�䂧��@������U���vU������ �T#K@f�㯁����|95<@���+�-�)�����K���FI�k���*@�m&���
���ma1[�2�u�I�\�U�yu���o�|��2����;�W�W�}P�K>%5�'�8���׫=����k��,�t�M�0�8]q3���Nܺ�^�5Xz��t�l���&��v��
.|���A�vP�}Z:�/��
�:nr��qRyA�}�m�V �k�Ш�u��F8t��f� @�����}��
�0���7m��*E W�<L}�c�N�l'����e� �W�g���y��]t����i��t��e�!a������u�ȑ:��"ī��<��Hl�����to��ߩ���U�\����Ы5 !Z�S���ҩ�ֿ �J	1�X�A�t]�U)?'{y���#6Q�K�ZCt�Ŵ����k���$}��V��$�_�F�CĠ�vbm���ˮoGb���ł_N�ʻ>f����A:OX͓֜��[�w�k}!�3�:��:�W�H���ZǺ�.�1���3���q��Z��D��6{=�~�,�����!i�L�q��ȽQ�l�d����U�T��&1��Ǻ1���1C���^|y*��]�V�;?��<ڗ-y�cE��:��E_�r��j�K�y,rrI��;��FAj��Y�F�$�X��ms�d�&��n���c�E,K�H��O��3�_�ǡ�}��C/4��� �V|�O��c�J�u:�z	]�*"���ࣉ���M���o�k���� >Y�=3�=�y��-Ltyq]�2�Zb��HK���z]<�TЙ ����[�����w�v��"c�H��;Sy�P�� �YD�I���4�V�����P4q�CIUL4+&MJh�-���V��Lq�˗���H�÷�r���������9*�6mv�;�p��NI��|�p��nEf��ե�{A(�O�P���x�e�a�C��˃�6V���<������Z���mj��z�t����VS��e��5���"pT�'>f<�6��̓���s�(	)�]�_B$����)b8�TW~��0�T�Zduݝ˵�SI B�vC��(�{�om>j"Z��A��O��D+h�)�F��V1:3��}�ݟJ%�l+�f�f9�"VRp��o�6c�2���3/����� <��}�e�i���r��Dh~�f�L7�tS�A�<,+=�:!F���蜫����n���5��x�������N���?Sy�J��]���㧀�P0x����ǫQn5��/$��P#\I��Mo�U�R��b��[�*��%n!�'؏�F�hR�`��g~P�Ed
y,��_Nj��z�ls4ejKR�S!E<܄,n�.�0�Ex�q6k��qF��Sԟ�`�Ԥ䙓C��YM�r�� ��%���-�9-��\�[TI�{�1+���6�=�<�	v���is�z�GAMZ�U����.<4�3��(UJ��RnLzYد ݂P�tų���I�-n-�Jf4E�]b�Qo#��l&yq��EwD��@����o�֡P�J��3#��qI�y���k/���TŎ�c�x�	���ϥ�=E9�(���>��ө;���%^gM��g,�����;ށ��*�A�0R}�:1������5u�ʵQ�g��B(4=�����B�>P�F1\�>��s��^��5�'��_�K���E�hn�ζ1�xŰ_��3خ-���^�69y+h���@�����V�k'{�{J��m Y���R,�)։t��:�@�Æqjk�����W����Dz�9�:��� p�q@�$�@%�H�¾~d����c�6sSHw{Ӣ2&�?�e�<�*�]�=�.s4����R� 6/Ң��h�|,��#�b�K����-� �M�&]���}H�k���5Yl>�'�<� �xݟ�}C7�����+��T����ka2<�9l>ۿ���u}F�����l�ZG2/�"c\�O�\���#��Wg���?�ӿ�(��h�!�ߔ������Оы��z�i��fp�P��d�R���L@���m<�HF�J�`�P��s������H�VX����H����{nx��M63����&��{5zǢ�$ �N��U���2[��32�w1���z��̺�p្6B.k����@���6�{�s�X%t�]S��<,CD�XA;Ƃ
#[��	 ���1�v�[Ea���� �`%���s^O�v&�JOg]�?�EAJHg�+LzNj�\�.�1�;�!�ÎbqX�X�=�?4��	�����*��=#k�l�0$Ɨ����y��aX�ł�ى!��w�b*�k勤˳恧T6���q��_z���	�yh�ܩ�D gj{W4�K,��>F�u�I�AG�2�z��5@�dF/'�ĆCѿ9��Ӏ�� ���z��b�dAY��m��W��2�x>s�r�f��e��O�=����3�F�#�  [ c
RS�]5K�3D�;�/�0鱑9���sE�f9�>}�t#��}����+�.W�4V�t̪��ɮEv$�+�˛0���h��˙tR�U������
��6�E$�Obfj괺wf���̄_a($CX�QveF鑎~G&g���m.|f�W8���.%V7V����]
\����ThO�1�Ƥ� *��l�/w#$��rɇ,���Pg?/c�I�r�	' J�/�$��Zc1@���&)�H���_d՛h�Ϛu�����r�5���+�$$˼ۂ(4ߡ�j�U#<<X��޵�[l	���t<&@�%ww��riU`,��/'�\��ܼ��턺�!	x�T��:���kkI���_�p�;���M�7EO���_��b�e_iY�d���9�\� �]j��mEF4d5$����Y�������.��_�������6
>C����j��`�J�)uc�
  dlI�|A�3i���к�.'$�\N� ���M��vưUS�0=�K�+`g�Bړ"��	5cA�|���"����LP=F�1��Q���J��.���Sҏ��'�&�ץv��^y��|�O��{	�}�=u�~:<k⬚@�]d�D���&�����J+4����g�.[���W�Q�A�鉵�����D��WԖ�6���H�CxE��G�Oq��X���9��&�f��FbQ�?A|�=�75oΪ\t�1�{{��W���c:�|�u�q��ɧ�smI�LF���tO�KD�+�9�!���֧�,���.��#�%��Ű��\�\���U�B�RX��������~z�p�\x�$*�3�\��&\ �h84I��b�艀����v�׃ ���}�Eܥ��*~�
,	lz�o��>������2/�BZ�9���Ks7�m	~{;���K2ɵ���3o�b�\`{��g���m�J�^����m���Կ[�/,���!m�^Iq)�����=X#��U3�VdBK_����p�?�&��[�lM�(�@� ��-�B�ljP2�ԅ�����U�
(�,`;�%�<Ty,:�5������;η�q��8|�Z��D�ePT�S�J�cV*�V:)�s�Q�����.�>��}B���-���Ն␸vzӽ;����ǿ�vI���>�ZqF�Adz5|j����|x��ѠB���`1�0�a��������v������2��Iw<ﬤeںr�5`���g ��"��L���ͤ�]���
vaE����k�墝����{uӻ\��Q�nl��s5i�X����L��8v*����q���N=~����P 6m�Q�bX+��>�}x�Ջ]�j8���G�Ǖ΋���m�Fuy��]�{�����Y��%�b���\P���)P��"����g���:}�wN�M��\i��<0]c��%B%���s	����ۃ�{H����_��A�C�sB��Y�T�)V��%;=��۴�8��lH���ar.��(�tХO�K��ɭ�L���a
xI�\��#?:�ڙ+�>Dx5iE �䊐���2)�� �9�|���E*�`�3��ݭ�1�hz&���ؼ��q��	�4���H��6�c#R/�� p|l�뻏�Y��׸;�W�d��>�c��Q+�U$�~�s��9Tը_/=�v����_~U0�ceު��4�ЅԪ4ӹ�ۗ���?�Y?L��d�ɖ��Loh�M�.e9<g^���[�Řv���w��2m��C�0Nmd q�=L*8{�������2�=OT3IO�������޷,\�ݟ=f{X��.T_C��h���b�sIq�;C�k1���1$Ky�/[N�I��?z�V��`�l��װh��9��Pل�L��=Ƌ�3	ܸ�G���o��sOV�)꾠U��fB�)'Y�\mɰs�v7���,p�*c{GwhJ(�_��}۔ް�-c�u�lE���b��m(�(�Y� �Il��Bя���l�.���J�l�~k�|D���I^��*@�����|�O#�i�F<����J�I�V���7�͸��硱��_hlQio�z;�Qe�Ob�ɕ��U�)�c�F��k��x���-wo����xy��,�����4�qP�3ɤpC���W�v;��o}�o�>}�Qh25&d �jﰺrkW�eŌ���eA=�@h�Q�3������[���1�M�I�lF��V��z�?S���PM�ʆ�'0���E�Ha��v�\�V��}{iU�Ǝf�v�{�T�ܼ�]��]�bN�̽��Q��Fl|8�#o+`ZOQ�M��=O$|;_aS_:Ji6቎O��S����<z2��%{�%�+Ȉc�xk�m}����������I�cFo�P�3�  ��1+Fa����h}�U�wG��(Ϳ�H�E�z���df�w����^�=3��B	�]�y/�P���b����KH7[7�g���?�����[��	��d�����,���W�I�bO��~��N��Υ�q�K�k2$
��=�D�I�Ck1����+���I*���Q�L�f�������ɯ���z��2���ר^`��� ,��Z�wTP��s!�঎� [��> ڂ�A�(���;������l�E�9��\r�UA��NRG�Uwތ���)5�����_3� ������a�\p#L�s�����/�B�ЈpyPi-P�����.�}7y��=�� 寐6�e���������m�{]�P��H# ^�d�>�M�y�D���� ��/�I.��WqS�f�����\��.ᆶ�K6
P����v�~�Y;25��]T�b���t������5�$��!`F�n���;����]�;�"D��ƣ�/��d��|�bA�a�:hs�^���l1k�5�so�%줱w�z&�٦
3�0�M9^[�����%��l��8�0���t�-���2�NC�b$@�t_	ܠE�Y<�̕/�hM��FQ�a�\�h�p�n�����]��}�$�����V�P�(���v�K�R�6���}��zۍ�G+�<;���w����G���-r+JL8y+3���{n�P `ۼ��&��VZ
�ېyc��Ψ��
���#F��eI�I�ȟ���	��槤[J�2I��_�/����i��mx��f�|�����J9�e�ɿ��?MT./u;V/�	�������!ݷ� E���f�	u�Xg��S��5b�ǣL��=+��p=z�*�
��kÜ��6����,`6%��W7�Ei���,��f�ߨ�준�� �.c����hX�����=\잼�F	дC���Z&��G m�����3g��5g�lQ`[l��5����7�F\�{�ҚC�l�U��Ysvm$�r��8�Ӫ�ua�H��[��x��+a�)�>;�A$�(?El�]�%ڍ��e���	ףg�/�Y���}~>BZb@�r��`��[׾��n�@sd�
�`rPwNr?]����Z���f��/!��l� �j6�f"	����VX��{�v��>�`�լ�����!��O�
��PC�(g?��\тF�˄nm`�ܧ+��E�\pN`�U�ʟ5be�d3͇������?��\e ��C��@]Z���S˕5��/e��A�CAǧ�Nct����G�zx�9�[ŏ4Rc��VǗڊm���S6���!�4 ���ݓ4��T]<���!�6m�9[�]�z;�ú�$f���#P���_�b���4 ;�4���Z�R�,/�������f+��-Y�Q}�� �E��@�Z�Ө��ф��Зt�<N�6���_C�L�x
p��`L�L���,�z��"�,���������_�������yR�6>�V`�O�V��>
��H6��W��s�n+¯���_A9Îm�[,���#N��^s��fY���x|/"B��\J����>0��Hhe{/��P�oq�Ê�@P�u��� �J��Am|c��a[�ܜ�yJ�4Yj�G$�@t֚�'0��0�����ص��d�e� Vi�9���RuW"�=;���G���T�:=�ʶ�|�zBx=�o\
��A��T�Nf�&M�5��OaV�=��iwBU�a��~�wN{�1��M����0B�f�Cff�y���lf�����?1�7~��&b���q��`���YY_���Zi�^�����uq��#eI��5�e(����ht�9�z����
i��8�ܸ
��BҀe%�3I~�'� ��0��D-k�4�/
)!<��0)�2_�ɋ+l9i�8�NO��_ ���d<���* E�`���[�m�B�!?o)�ǝO�6�b]��EqV��i�C~e���J�(�&~1�i>K�nt/�����@v3y�t}�_�D����+Cd�HK]^�_Ƒ��<D��(�@ff��/��x#/c�\�jӄqQ1"s��=}
2�o�!��o�#���؅�O�f�sq?T���OC� �c�*E5kʣ��0��8����� 1�h�*�^��xӻ��"�c:�(~���z9�ӐTx4iZ�&�M��K{���W��«�I����5���`Ԧ)\p�Nyx�w��̵ܵL���|���c�݈?���`�f���Bp͌���7!P<��� Ϩ������J"��7�Ѩ[$<�t���]S��:�SX�1��'�Ɣ]��}���bt��E�2�3�~��=O65o'��H�%q�t��{��Y[�Ӵ��0Ph�)�y�)�#Fp�e_�lt�vG#�ϖ�w�=�xn	�WX`	��#�$���x�L�Z�BM���]�l��*�{tu��׸��AB���	'��i�rrH���;�������x�S�wt�\����(���}�"�wD4������y�8;�;���J���[7a�0}N��^h��[D�B�46��%��m�֩���;\��y�8���Ѐ�J��v䂖)J�~y�n�F
����~����x� %Elr�9ỽjς}\�7��e�EL��{�$�{ۅ�j��\�q{�^1;�)0���*jv��'G�@ ��55o��.��������2��kЃ��?��o�D��1̋9��TQ�G�ۛ�>��[]^�F�e!�v��mVc:6�4���Z��O�p+%W��N���xe�L� �r����?h�0���m�g�R��Fh��fy2��s�_�W��2�*0��z ᡰ���3�7B���@p�m`����ϕ9�I,��Ӳ�3��ȝ:�<�oغ�D���5��;�P	�J@p����=���j{.�9i՞t.� tСJ�Gۼ~
lL�<��`}44>��D+�9\"�r�eՎ�m(A}b��Y�2�#`A��p��q&Z�W!8j�WC�x�e�z�2H:�e�!c��mp򕘎z>��@|p?���m��lN@mK��>��6d�*�n1I��5�p��YN��m�7��c�UR&#-��֖�-�U�����B�̖��9��⭼C�Y��& �~���$ǲ�a�L*R���ai������a~&#zN��.���l�6�H��ڳp)W�z�w}�Q���\�U���Zw���d��P�8���FW�燧
0�I��כQe�l�RM+�t���,;"�>F�"��=�}�י7�?+�]�yP_�R7�5_@�͸q��+���5�5��q,8/X���W�P\
��� -uik^w�sҌrMf�)��g�p_6<:��!:mw�_h��:���t�q��J0�<�Yc�N4D�r,/�m�����?	'���p� ��R���������huU�c �Y(�� >`:�~0ɀ�i'���w;������Y�A�GHD4O�l�����,#��~�YR�cuh&ǲ�����6H��D�g��,��ւd�{7�l���8�����xq� ��1�k9ҭ�>H�ז\�|����7�AD��`*2����XC��zG}�=9sno�;[�iN�P���^_s���<7���cVѤ.T�aZ���X�N�_TإZU�Pi����!����<�n� ��-.�JD+��{�s���=�����Lk�*%��9�W�U��-8ٹ.Y���;�=��5Ki�r%v#��18q��+-���W�X��,h(�E�ѓ��Y^{�]b����3���/��Dp�:+��S�]['�`���{Z_��o���Q{�tE��@��-"�k�ؤq�H�^ !,�
�z�B�i1��W��m~�Wgi�w-K&&���^[V �<����=��"�$|sf�:| 0��ר!UpR�f�;}6���P���[���e5��J-�^���7�{��[ܵy�f��C��_z �E�{2�������6�����լȀ"�������Vq��f-R,��/�j�@b�ǹ#q���
P-�� %���Q����]�(C��)�Ϫ��ž�������i_����Z�����u
0�I¿�������^j�~q��T����� �=�L_%�˽�X��k������6yM�Z�*�.���/k�T_˷��� ����B�e(��$ĉ���xbZiZ�Cqƙ���K�~���8��� ���t�a��释\��G#�7���]�z�: �m���|��&p��I)k����P�(Z��΅�D��������
��Rs��np�Y�hh�rUε-�{B�,zhO��}h�0�U�b�A��c�5�.p�f�ٽ!�@�7ivL�,]9)���.x��O�ݽ�h4��W��C�U/�TՎ���'>d�ƾ]Oi���%E�j�.�,lx' B?�Ŏ�4�m��'���W���Ynå�9���(_��ޅ�GS�y�f��];{z*q��ܯ�mP�d�(%��T#�����g�Z˱�#�zfg_=���c��\G�T���r�k �c�^�����1I󗪷?��أ�:F@���V��hv#��!�I�D�[��Lu�,�cSN�7<�~I����Xl46�д���2+�K�>���wVt[h<˜��M�1(A-��n�G1؉J]���/�3�,B$߁t���Ͻ����H��{X-v0�K�$��H�m�>�W��I>~-�m;\�"������p�-�e�p���D �g�����[�/w��.;���8�D�ы�31�b��QXbx>nSU��~�����7rV�{ ﱠ�q�fj�~��ο
l��5H���wr��C=�����v.C/���9����У�:3Ҽ��A��|���e���1�l�pv@�c^�А�'g]��,rP�kdaM�5�K�ڄȅH�N*R�wۭj���w��� l���LBX�·�罧�*b
^Ʉ��1:囸��a�*cZ����|� e[�Jh��5$��(�0t�2���� �g��9�y=W@�I�-�r�n��e	bO��t��:�ɮ�n�*�&P͌���Oˏ��
6��i�<K�I�c?�o�?Z�������lEL�L5����������Wl�"c�NO{�ni��� ��k����2E�g��Vw�)��`�ߏZ0�3��	\�xu�d�SH�ϑ��t��M�3e���2~�����1e��1B�s�q�`r+�0�%(�m����%�MTo��T's��E�R`����c���fD�I��~92�L$ގ���O�mC5�Jt�u�4���Q���z��7*�~�����`ҮN�n��lܘM<� �ڜ�ݶ�*�
/	�ou��WPa�<k|M=1���-˾���(F���� �B�6�#��"��S5K$�v�ʹ(P�y�z��"e6��N�P��\!7Ȫ.j�>j�&$x .+�-�>���/���u��2�a?F��!�4+�&����|Lt|¶*��8��y�{���w�@Xb�X�x��T�5֮��y���OT���B@���+�����H�`ƹ�g���"Eǹ�R|�í�V`��X{��4�5P��3m�㰥C(1�Am�!ѓ1���m�"]ѻ�~���.�Ӗu�+՟X����EGG/"\6 ���Ғ�:X��#ݏ���N(UM�)�Vm!,����Oa Izgk޷�T{s���?����*��e�����-�r�F���L��n�Òue���p$�����3�(��܀0���a�z3��lӑ��6�X]���)u�.4�T�)�w��G&�u�e��=��S.M G�)
�A�2#�w�U���./E���v ��y�ˋֲ�g�dXӀ�_�z(�"s�	��̐�����f��\
`qFh�Ё#�Zl�^� �ơ0~O#�w��t�)��bDcTB���e�� �@�^����[��Hw@J]�S.T9��_=�&�o	�H6lT�9����P�СJo�V#}Gj�<rCd+��\oR�Z.�[���|y?�����b�
 �"�
QL�<�� b�1�kI��Ҳ	A'��Z�ޒ��*W�L)"�!�yYN�wf�QFte�\�[e�����|\�@T��k���&gv8��YVy��)�[�(�S񄀼'y.��d��!R��#뉫��H�X��[�Jl��u �D��=qh9M�����֤"�:s캼�Wx�-K��j�ɚX�/���GS�sE:�'\/�i�� �����1-q<��=(d�e�["K�3O%#�ķm��4;vWJ����ڗ�O4���|�c���cʘ�2`LZ�y0jV�;�
����uU0�&RBʭ���H[c�s�)��F���0wP�O4�IŲ��)���?�9s�_q�r��d��(����4��Aum��:z#0�Ԏ4�t��3��Q���O�YR0����T����(�ɻkfM���!3��fWm�K�P�|�����I�'E��:tPP�\l)��9�)^?�'t>���=^!w9��m�/%F�=P�g�d����"�9�� ��
�V��b��u�츸l����Sv�:>gH\� u,6���,���v�O�چ ���t��v���.jg蹼*1��_˵�� �[��yZ���~�c�����(J)L�����L���E$y�%���Q��Q&��#�IO��n�nb�i����K��2��^ۙ��?�i�"ѐ�ƿ"�6}7}��Jx�{x	��_�bw�����fhpdÌƗ�����'���B9�A���.����蒀}k? ��R�VpL�N!S ��r��:S���9x7�֊-� ��&��8��V���P���R�(�&:�}�Q3���<n�:��յw���w�:��YdU������=/��颔�����R��τyU�i@�R���;m@�Y]<u��=�&J�-@�ʋH�~"|;n����]G��&ʦt*˫��w���a�b�Um� ������o,KƊ��`1����!CB׈x��?\���q����,]	y#����U|������ ��U�$5���a��9��0`�<Y�5���er�O[_��R�e�e��/,�
���?��\�xqs�	z�񒼔����ݛU��[����3ލ"�.U�\��Gy6]%z��h�/�Ǿ͑xo/�ro?��cɃ���`��Wk����ز$���_��9���XV�pv4��#�Nt��&.�if*華M�ʬ1x(��#a��ߨ����L*�Ckb��%0���YW�.j�]ˁpYxK�\��9�VU�L<�!S�ń���N̄�ҏ�&��:J@
�^��z�|�F${�ؕ�i 74ׄ.T�Y~���x�	W���>� ��A�y�C6�[�s�����:U#���Ľ�LQB�<����K�$�g���#d�]�޺���$:aᕖ������>��%�W���+�.l��Q�D+�O-�M�(�݌�a���a��9�K��N��&�V�cg.���Y�9��F1�#H�Ne}�����G�70C�#�)P��ZÁ�y��K�XO�:.��i���ʎ��@�vv���3��z Lp)�|�[q��HG���D�g>k؞ɜ��:�4%�i]���]6����"0m�,n�,�m�{f�.Eu言��,4$9xw�! q�-LRw0���-�PƞVYn�Y��(�����0���|� ��?`��*���-T=��8�u~�Go�T�Q�=�>;�������3��Eх���
�la��1n��1"����L������]k�����3���;i��B��#בv��0������c�CM�yMWz(t5��ߓY�ف��O�16)	��)K�=R0Y!��v���g4��6�Y�
s�C�`h���v���"B�H�YF�=��˂z;��U����q��䅓�0y�%˥o�R����l�-k���_ �O�G�?�y� #��S�`s���K�lE�O��M�lc�;A���`ajA� _�\���R,���̓����95e���iT�U��-���u�3�r���}�`�n�!+-$!M�-[�f�#:�O�����Y� �~�*��Fc�횱}��9�q�fѾ�J���iV�ƈO=b�;�Z5��Y�l�/���+�ק��a)K��{(9^��]�.��_�®2;������E�� �^��nc�p>/[�U�XEj��b�L�S!�w��}S�yl��9�Z�,��*����,�u���g��A `�0�$u�U�hJ�\}7�	SLݱ��K3+����u��G}�4�h3S�X.xC�(���1i �o�(�F��\�E��¬v��yfK�$��.���ښ�A�I�Kv3����)*���xIЩw|�TM�"�p7�\YJ��g�맔�g���^��j�l1�[bF�^~S�1c�ĮP��@F���M�ҝ� <~��
��Pج-���.3g�n�o�sT2^�Vpz��1`%�֎B&��?��>A<�c-�K-�&)���̽�lv�H���z�X.�����t���!f���N����m���E1Qx���ܑY8�wɠ)ABP�Q�����ꃽ�i�#���׺t�z�\���ڡ-����yW��71��^��AH�r�](WN����L�7aƖ�4!��cRQ��6�H��s��̼$|1W�E�57�M��Z����n�v��E��� ,#0���9連���][~���`��_c>��nY�}��o�$�7�9�!��LއV3Z����],����Y+�H8��'X/+� l�W�Ct\e
έ}��ZZ�7���h��A
�o_�hԴtb~�8_@��nL?�U�-\�?`�B�'���z���6ݶX�C>3`��#�2�|}�G��:�ċ�5����g&�O�4�I����A�L6+��$Ɯ��[£�s�~��U��٣�䶦��W$�je6#{w��FP��P�l<��������}��'��A���Z�V����r)�%\^x2��|^�H��0�Y��+C�T��M/U��#Z�Q%�IA�^&�����g��E�;�.��k�y�pR	=� ĩf������Ԋ�9�ͭ6��5ԢwFR-��w���rwk���l?�.��URd�L��#�p-�s�g�������>"���`��}��;F5���=a�{���ڒm]=�B�4S�1�wS�z��.��/�ʴ��0��5�?`��
n�b��-�ު ��U(/��$,u�&ޥ��XM�)ҿ����B|)�j뇮Uu�s�N,�IT��!��f��\�|��gV5�s\�6b���%�z6;�U�����q���7����螦�	��C�ϖPX��̊�_CP��kK���5����Ys��vX7j��V��:8�z`>
)�ǂFR8[S�oN�wjV�./��?]O�p�𮳷�_\~6ͮ�l(��x��>Y�L����=���)U��;��Ǣ@ڦs�]L伱Wx2����9�Uf�IH; m.��i���M�Z�/��SO�� ?e�������,��מ-���� /��4�PAF�3R��$4C�`;�����_:X���Qfge�_����a)��͡���'��ͅ��Y�);�]N�vh�H��D�� ���s�!�mՎ�2+�����a���#޴����2��3Nn&�:��|�������	��d�XMU��l�LWé -瓊����D���F�^S�f��<׭w���w���|�y{�Fr �a� p�j4ɹ�9j��{�]x˺ P`�8����p���-E��1W0r��-�JBb���$b�\�;�Ӈ���S����L���g�����^[g$2G�����a�嘹�(r�*|���,�x���+�l}�1ߑ���	����*w��Ɂ�� a�~��=N�3�x4= �͉��z+;�x %�r����>�`o}����1X�
GW��ɟ����Ǜ�sKg��TT|�)^j��eʰ�r�sd��ό�s��`&�����l�mIȭ4�s�J��K|Ff�: E�ņ�⩓4�K�R�ؠ�1�I�����c o�y�d�[�IC��X�M<ƶ_��+:�^�e�W�+�������A�C��T�f��^QK�R�]]z@�b�27+w�VT�W?��=VN�*8
�͂&�I�EN��"�������-d�<��^�ˤ(�hVt������OV{�û$q���zr�PZ��Ղ%N	���r"
6�д[�>iM$�������@>�^���~�U�w!#S�� ���^��/��{8zP'�AJ�R�٭�+�E�d^�?_�������\
w���8����Id�67��J��f:���oq�}.qސpElqTi�����u%LO!&z�{#n��s?�;d7�v.������/`P	�bE��T���(�ryФ},��j�6�l]S^�(~��N���(���(��.iD%6=�*��ˋ�W�V#Տh��f��	ؚ���gS�h* dv)���F�W��_���yg8|�|/�2���&�6���ì���*�89�@M�<c�Q�C�Ayw�rBY��L}|�n�i��, ���i�Ɲs�}@�h2��RųbvI�M<>VDIߢ�@�����}ph;������lh�4� 	��q�X�9���	�;$8��*�$��5� ����l�v+ؓT�l(1|�)V�P0�'�l�vRS����}W,fL-|��|*�ډ�8EfE�u����N�Bظz��������b���BM	�����a\�8Wp55G�)`0Ӂ���?!G�%n�,���t�vf��t��٤=���Ӆ�ԁõՎf�8�yw�M���ۀK�p�	W��Z@mv[[l�Sf�Ad����(bo���O���z���e�j��[�q_,^���u�@���;�uN�Mk>��)�M�pp���qS'��|�"֎.����/�� ��h>K�x�G�_;�