��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$��7�4��L+Q���+2�"H�������v�ao4��	�u��=��d=�>�iV�f��l0�Zs��7���~rM��U�`���e����K%�u��ݒ-� rā�SZ )����C.��&0C]�-��[�3�-���+��պݣ�k�J�vo`�A�����f����u�X���v�=�а���]Q�Wۿ�߸�=_Q�X����j>��Zw�K��SvX��ƥ.���#�����Z�0���#7{��\S$��@1I�QX~TQ�E��db����۰� ���>0�%�9�j汈��}��1� ��2���h�G��SeY�a���	'<x�p��k�H`�H�j^y�0�s�78+���ֳ�`�R3dW��_��{p[�?$�s0��#�zS�_��bH
�c�p�IL7]� |����Q�� ��Rr���=��E즕2%�����`�^��l�q-�]�p��jf��Ӽ-f%H���ȳ�>��+���M�71��4_�) 3�46h�rb�J�W� k�h~K0�>P$�_n)���5�r�j��W�J&޴o��$>��6��ŀ�;A~<6P��K�~��f��*I
�Z��}`q���ApC��n���g���3��-�іrO�mF���,�$��@�BI�q�}��Ȥ֐����î�䂧��@������U���vU������ �T#K@f�㯁����|95<@���+�-�)�����K���FI�k���*@�m&���
���ma1[�2�u�I�\�U�yu���o�|��2����;�W�W�}P�K>%5�'�8���׫=����k��,�t�M�0�8]q3���N���GvZ�i�+ C�e
��Ќ�S�v<%���q��e_��
�k�夞��>ZO7E~��5k�TW Aod��eE���G���ɑ-'���?�G$����ќ����8ɸ+ 5ʗ���l�d��,�J�
�^�3b,�����J����#n�zK����z�&��;|�\�^���'e�W�����">�w*<���=�O�V������0g�R��6��X�CT,�%,4.�H%�~�׾��-��CD��G$���4J���+&]qߤ�3L�T�R(�Ӌ	���!>M(����m2�aw�H�Yl��amE��V��r�b:��nS��Z����(b��>��Ͼ_V���!,X���fQt�(�kQV$�7X=#��'Ǜ�Bg�K�ߪ�� �����A(D��)�,(�K��^p��3����J�ΰM�ٞ�}���j^��B3���ǧI\�a��Q�qn}Sd"��u����}��[�ލ*�6�g��^A�V�C�K�GH`�{�T�~D9�@˂34�g�NF#J�����I��NyI;y�a5���ؒ� ,�?����j[+�R�KA �^-��W`q"y�=�'�X��$�O���Aa%���ϝvl;���kȜ�~W����1�tΒV��P������!�Z~�V�݄�#��Ho���]%�¯*EiU���9Їn�Hՠ�gf����Y�邌���r� �u#z�!�I����3T$^\�T}�{���Я5��gd>�΍N���W�U��������K�����]z���9�������E?����d�"�r�={)@���]������nCV	K�@��˽O������(o*��5�z��i�q�vs�+���5:��'�_�����NSCI����Gj��=�7��'%y�X�|��w����8A�=�,��B�*��$u_5������e�-F���Ѓ�\qѾMJMwn�u�;d+2&z��D�d�oQGeO�0��pr�<��l�#Et��y�t����*��D�I���Φ�~/�]�J�ؤ"���sa{�����ʡ�ʌŘ;��w���p��*^�O�0]����c�Ӷ`��\&N2�K7 Q8�A�d�Ϻ`_t��p<.��_�FD�k4jL*2��s
��G�m�a���EH�(�^U�%$�U�X��������`7S��7O�U�t�/��8�Y#�Im`.�^���'�&#^�d-v�o`��Ƙ�d�Ϙ%�Y��T�3��"1�^ �2�}�~OK�c+Oy�8���:�dU��e� 4ZU�V`�)��C�:��1qn��ZN6�m�MC�xid�g����C]V7� f��m�N�w��(șՈ����"fľ�^%D�#|1�(\�~���Ȟ�vPU���W�T@BX_L�Ec>����Y�p��K\>9g�U�Lñ��F ��ڱ�d�sk�畎b֞?�	�$S�A�a�`c��Gm�,@���@�F���r}�ט~�>\�\����lq�n�/+��E�z��/[�f�}Ɠ�ך�V���o�۟tn�8�7<K����n�n��*(J��Y���T�:����7u���R�Lj���t�w��c���'xƟ�*��]|eI)�����躃>��9yi%E����q ɳ��D}Ҷ�"/��tU�BS��]5I��z'j��1�77xc���+f�n�B��ø��U(�] �â/f�-.TK��%�~\䀘�lL6�"�[�L{��ȭ]
��Z4a3�f��#o�j�W���S�
�{���cv��`����-0�}$pH-�ʃ`�-&��vG�6�Т5��z����B;�|����G4銆�3���\M�����ٟ�hNM��LٚQr�q����' Z!�Z�}�z��g��X����	 ��'H<�#�]+����)�.I�x��z�^���[V���
�Ϥ-(S�����Y���,��g��)~[�d��N�34ە���Q	�-���޿-d�?�ls!���#ߤb�H��Z��E���\�k	�W���C��HΚ̲6j-�#�6�X��e
��@��`�/�I�̪��Q�M�oW6UK:b(DI~�4A<�$�z���ۂ�D�{�y��5v	e��� �WH��ݍ߂�#��M�6�4	��<���|vݫ�{�����$Ww��q��ȓ�9�ca��Ga[��ױ �$͂g�ݫ������̺W�����tH�0���%�e`8�CQW[�p��p�pnS�l)��W�.�	R��<�	}J�i�fb7��nh�l5��Bʞs�[��[�����)m� �����yH<��-,_S��U�ȇS��!��Zo|�����4G���L?wK�U��
.[�uΒ��X�S��%���j-5�&D��
aT�N��Cg��ӧi5jR:�6i�^��D፾J;�OIA� ���`@�:��=$g&m�T>���&�X*�˭r��K2�j[�N�:EߝF���ű(��%���^��"�7��$aw����ntk����f�8��y{�������.t���uv;_~ q^�=O���o��҇�?U�5�T������4G���Zc����o�K� ����
����F�F�
����P�p��G���j��C��W$�	��3U�GQ����l�}��S����D�M����A>,�ʥ/�o=�J���l�b���;�u��i[r�4z@���ށ���If�ߠ���S�|J� ��@+sC�:�O4����ܡ'�����r/W�;��̷�i�� +�7H�,����k5v�|���j�-[�:^k��!$��{I�($����*>�j�z��ş(��0Q
��ʟ
����aW��vr��&�qޡ�=ye�P�Rv�&"�����z���ۉ�jJ�,��{>��F"&�GM�%��4���N�Y�Ҽqs�ۗJ�-���ɘ%������|k+z97b!����!��:�2�Y�Iz@A�����044&s�ҏ���M������N�r�o:o�}Ўb����f9�֢.��&}��~��ؐo�6/E�/�\��C���Ԕ=��a�XJp$���2��A�Sz)V�R���3��+=H���
�uaV��7,��!�{�HJ�d������z>غ��QV����9�N/(�v-,q����^�R�j��a��	
4��M�����R4�J��&V7�)����x壶�
7釁gUG�g)����"�:v7X�������F(ʘ=��w�t����a[W������nd�?&��pa���ٿ?�˃�I�|�\�M�������?"�o���Um��ƛ�e��!��zi	7���H�$����_�,<�{������M�$V���P�,��y,�hn���5���6��H�1�3�R�W�T~�wFd��BH�٪y;��B��6�Ճ}����Au�G>��{݅UǄtY^��G��	M!Z�4�=Ь�"2�46N�5��k�اŭ�[��x�,��6k)�θ�E��oIͮgX��1��"2����;[{N8ES����a�^P���<�Y�q�XZ�i̮��+0���~�4س���t@8�gD�;���4)T��,g�?!v�8�^��f�X�h�`�q%�yG��
��C������b���j�Ǿ4�o^��pe"�a�*�<а���:ʸ'�}����&w-���[<NW`��F��A�N8]\(g��[���?g_01eDC~�|��}����u:�*5������M��#`��5���%h�C�V�d:3qY��k�.Oo\Y��@xp蠷*����r)�Q���9����G6��zpG':����IZ��{_Q� �J������AQ�L�(�r��:�)r��'��wC!��s�-�Xt�r�\�w
QI?��ܢmRd�$�J6�0�1�*�����{���|�	���f��f��1
Y�R�^aSƗ7w�N��0�԰�����Y��8�6����SZu����n����0Rm��ȴ-�<�zy��;F�s̭6=&��PqK/M>��
���9Z����u�2�Y�k� ;�13�`Po�����%V���G��U]wS�H�b<Vo�>�NW�b�!�c�����]u��R���ҡ�63�{F�g*��~ܺ���3"Ǔ�, tX�h�p�XM�Zw|���������B��՛�e���7�D8�C��I�3�Z3�Q�c��"nҩxܺ��g���%���9��B<��<�ȡ�CQ�]i(䒁�~�֥�)aG���v�e�{�s����q�W�G�sǠ#�R?� ��xݎz�@�s�S����7?�bK��b6�[�pC����ӋV���50���ښE%$�	��~� F�J�I����絳�Ec}~��+�y\��@v�7�w�)0!y���%0���,��hd?���Z�x�R��`��W�\f��}@��S~��`����7`D�wd�8+�﹯[,���w��|0F1�ù4�ǾHS36�ў�"��KY�4[Y}�H�����S�3�Ki� �72���Y�qё�f~_�f2��ɡ�t�j ���O�_7/�w�9C�4@=nhy߆��Y�T�b^F�蚢���p�ޒ�嚹h�W�7F84�6��q�)J#��5�ӥ�90��:*8�?����=�����ퟢ�ڰ��3��/�k�BSq��?&�#�,S�_�1-68e~�0k>�t��!-*��
�SlN+je��Mb4�jevC�����]╂�$6�L�>�2��x��D�~aZWz���ˊ��(�B��6�7�I�ܧw�����ׄ��zh/����I�d�9��v!'o��MN7�ߵxO6D끪h���2ps?��f���G�sD��`�Nv���Xk��1 ��9鱫�̢{�45BA�8>첓,Xdmݙ�S�f�J����*>]A�C���Lu����/P��'6'fύ����}C��O���R�\�Yg�_��\�8�L���O� V���k�~��R'�y@&��5^6�7��ޙ=)Bot��%����M�]繖N%fțt�����'�#'kE4�`t��A���`�}��>�]\#�g6�ft�ل^��e��?����������OJ)�D����f����fh�(<3&��Y��($���Vv)��\����ִ��9z�M�������r&�}�#�򢤓��d�ԧ�G5�t���G�?|���o�c������7 �:T&�Y7~�� ��h)�
ʘ�:��W�-I���Z?Ә��޷��g��>��W�c�4��1�D�W�0���\������������%�ٵ"�hu_o�y/{[4�ҳ�XD.Q��>|�c�a����s7<9W_bǎz�3�����g�����H;F�<�ݟ���ѳ����d����xo�烓���Sq2���%�<H�������ҽeF!R���A[���pc{I���L�	{���h�m5�B�e�c�<�0'��Z9U'��]P��I�\v�>����xk�ω7��k����Ι��� ̳u���D��wc�.L��Yv�!B+���G��S��ʕ�i_#���S���g�=��◨pjf32&B (q=��I�ib�.�id/�cqV4�:����U�o���$S��b`?��N���ޅjx[� ̉ �����i��-�$ ϔOS�g˻ӥ?ڵ��wxx�����z�OR7����[���^��̥HN}�"�� Q�)������{��X�˰k�/MM� �Z��xW���儮�#3p��)Jpg_��|X+��}N���f@���ˡ�XJK���￥s���"�hu����^�8ր�O:�JD�
�B�M��ʳ+���$�������,+���nv�HE��ܳr?�`E�G}�]��9�ы3��b�7AX�>�`�4������oUj���y�M�������^@�z=��*8�#�8x~�<@�!�m�4Z��ρ���^8S >jm&��6Eܢi��0g��/B%)�O%w���^�-f/Rז��g��5¤��#�N�������,�8�� J����#����)�|it�R�z��G�Rn
���{Y���
�j��ǖ�0/�ۮV���5>YR�^ =1����=b�����k0�̶�B8�f>��G��
��$�����'��j���a6�rA�,���ǵ4�
��(�gDCb�������|ZY��@�=�ন��w�x���-p���)G��6�D�5l?�?("��k�X�^}��NȺ��<&��e���Dy�S`OxL������gB�L� 1q,�>�j�a U�x�!�0
�	��ھ���A�ʦ[I>r�J��f�-)�6٣	8%��@d%��������jc]��;ӂ4���ϱ�T�� ��B��Y�1졅��y�o:�$�%5Ls^:AP���#oEP�,:\�?�M�Ec�վ�;�c�L�q�l�Ɔ�-�NX�>��4u�N��M�DѰ����c"HE�˂�V'�g��x�������Ēn����L���p�n3��J�@�/}e��X�F�*��j^�q`@ |O)�H&�;N�/�.j7����c�5�I�+�_cI1z��ʃ�)s�ob��u���|qD�������4o�k>>JH��G���= �
�"d��2l`�]�B�����E�v��8�
?m�
����6fi�\2����Ę�enJ�
����`^d���o�b�ʦV�}����#�V9��Ȑ���<7�F�=�$��߽��&��Zo��N��"���ZM�)"��<�;��F���[k����H~�]���=�5�BK�%ڢ��Mny<���b�p�ZY��s�
#����5R"����ظh��V���ܩ�b������S�1�Q�I�$wY�W���hp�8_3=�A���S�zȵ��
2�^,>3���Y�~��C���F����i6��0�	��C>�\=�v-�.�I�!8��lA����!�13h�@Ŷ���l.&��՛���2Mx55�/�*�\��C��n.8��F��Ln|�B�=+`+u &L~Kiէ��O����+2ó���?���@��Fc�4�s�{��f���?��h�m5�p`J,;O�~+����"f}S�f�O������/%e:ua3�I�P�*5 �̋f��.�$g|�:�,����sXL.�7f}���7@�;k��\��W�4�+[V�����AE��r8Ǿ2|6��I��M۪���倞�?;��ʪ]u�>�g#��m�8�^�{Ŏ��S�^cp �!Ha��=<�����1��b�-_ӡp�����o���;��S%��t��<���_J�>�%7>���b9����ԑ�"l��%�Kn�iIP�}ۑ�
�AU��Ҵ���0���+����;��sJ+���h �XeA�^��l�ѧE�f���>!�L�mȼ�t5�?��r���`<�Ya��p��;�pM�֜^;���)�1���"��hҁ1�*x_)��K�x�<�3����)���bdg����v���i�O�Kx�������̓�Ɓ�E�3[Ӧ�~�h|�|ú���2���C�HusE�$+B��Җn7�`��H�<�Wk*:�s��fJz������i��+섒W'(6 I]�ݴ7 LE�P�rꣷ�&��9��OS�g.7_��/�m�6��r��ƒ2�&=qʶ��¼����\�'�R�A�(����V�$��r��J�w��E��B"�^�w�(��!F��U,qO��d*����k�|��1���@�1C>/�<i��w�ί)<I����#�j��X�,f������e����iYbZ"�/*�nF��t/�ǰ��b���"]�V;��l�:�s~�'sI'WR*vS�t�P.r���i��	QdK���>�ab[�y�7,{=����F��cMdL7�(�i7�x1�p��:��}^��p�f��E��9C�~E.�?���߃�q�7�J�*]_o��zF�~����	�jvc�Nz7��$)W��Ue
u�r��7/_��՘9���Q�*H'�{'��3������ �����*Uj""_�v}�#���:���R�3Ӎ���C�o�k���U���vA&�2~F����[h״�V,���1�����$u
�V�����e�i���6UMw�^�%��%�K��������嵅���G2��2&`~�Dᴗ@#x�-�>tT�ي�A,Y���$�]j4�]�NTF3?l��$�==���
����m��T���o *�}tq��y���.Kq�k���<B�7�8R�f�ają��q[�Ѥ����p���.��)�Q�_Z?gv�� �
c>ʈ*�$RA>���u�.��������2:S)G7��){.:2I�B+* �6w�����&N~?n^�٭8��zb�:1�H��_�[������H���Fg����6�U���ׇ��E �/!�@�����z��d�f�{�����F���DL�Z
�פ� M���l��=|�`(�h@_�m��-ق!2ü3�2���蘩�q_e�['P�LvV���uA��r��@�R�t�������9��N��tE�l���\e!´�P��o'�҆���g�`/�J�/r_%n����b8\��g��
�p*�?���(�1i�O�*�3��uO�j��w�YD6��1^r�`!�� yl�����/��Sy��d�)U�j���	��r���ԋV|��f�J9Ow� ������0�J�.���_�v~�Y#���?��V�pv��	�K<��Jw/�8(�瀳y�>��$"E%�ٷ�0Yh�Tm�i\yW���:+l�/�y(�.� �^�ӄ���V(�*�Y�����qO�[~W#g�<-�VU��"7�4e�'�qI�{�u�<�*trV�/�����{��̯���������I`���~�Y��l[�~?�?��<�6����Ҳ�c���΅���b�م��	<���`�as �A�(@v�en��&)"g����[�b��&t����k%�v�������)�:���d3��Y-z��:�*c��Q�ᒾ	+�\im�l�2/� (�`�BvO���Ty~�>ĉ�d0fƴt��!J�9��|ü1�7|l0]��(��7Z��ĦakEh1���w�-������<�L����Xqߩo��i-V^U��6ތ�ٶ t޷��.����N�D}"w����PR���$��wC�!��G�'}Y�p#�DH�qfS�&�]�V��c+<𤶃b0�� ڛZ�EZkKli�`�����x����FY�(EPc?��f琂(��;��������Q�6ە;�LiH.d��!�ŝ�IQ[Iiܝq;_C2/r���PX9>������Y��t��23�ԫ-:��`�_�� 8�ع\�(���xi7<#��Z�&_`A��@qmϮW���L��D��ZS_0ԙ/�Rd'\Ҹ*�3+��6��(&1���P�K��:�΄����OP�0#c���$8�|��V�i�z��%���)d��ඌc:5~�����.��:��S$��?�uڙ9�\o)~-�����4��;k�2�ʱ!�$ �#?+���B�QU�m���Īo�u�5:=�𓶀M��;��߰M������Ci~�VR��6�ضQ-���j�(��Zv���p�坪�5u)�:�qAC��\�(v��8�@k$uQ��U����G��H�2�Ͷ��ǡ�j�����̺;<���#~��S��O���������V�䗢��/�h�CO����.t<�E�����3K��Fi8����Q��df�bb��>/�a�m{v՟��8}6���d��T�tW���C��eւ�����2Ā�=#��YQCN5u�#ͭ%R�rه��kW	���A���V�NK�!d|��]*:��I��|G�6��\x��D����~��G����1��joȽ:2�7_�*��)(s?����<c�P�� o�󉙑_E�����7İ����i��ou��!ќ���.g@�\g��wD5��k͕�C�/TKP�AT����/u�˓�~Jp`�ݢgv�����%���QR����ۮ1����6���������i
�=������DC��ry���ܻ��B�k��'��� �=Ri�{��4�������wct���|�Q�P��{ӝ?������o(�9*L�	�+|�����CW$GH7W�'V�A�[��ŷݎ� ���Fz.��r�:^�y�a$�4����HY�_�
�i5��!�s��B	!���%:t�C��Ab/%QM΢�|�Q�%�'ē�:�1��@4�$�	&�(���Ê�]W'atE��NI��������]�����92x����+��YP}'���Ab�9���=��,ӼD]�����C,1̂�A�,J�'���[�K%f����<��z̎�����JM	��K�v����>y�N���=��0&T[��I��1!�R�;S<N0;�
L
-+���H�sO�0n+G�'�������O��2��5�^�ʙ�pG<�ElN0lR�jW�1�7Gd���M��"|��4�qSg����4 ��^��$}��6ۘd�J��~�;R"�M�m��!�V �"�9�Áp���l뽸z�8v�p��'�j���	|�r�6���4��h�L��{T�ۡ��A<�{gE�������b�����F��||+Ɓ��SC攠����n������B����D��k�v�(2N���n��ʓ����꺡�k�i
��q�����_�6핛���`/��Y�!^vB�������3e�M�jƓ�"�D[�N�B�Ah#��PF ^���q.'}^A�^k'6�4��:N���A�F����0T��Y��:'���W{��+�;%J�/�o��~Đ{6m�F ���k�,����-~߼P<���k��M�4�u�m��dJ!�&��%W�$P��g���>�}�q����6��2,S�W?-Gk�Ӟ�*ɿ��Z:��mHQN
�e���%�s����z���qp�����Jt�>��Fk"<$��(ڿ��,SJ	 �w�x�ۗ:��c�Tqd�`��h�6n��ƒ�wV�b3P�2
�@�;ĸ{����'1��iWM8�#�Q���Լ����ĳC55H��k��rz9�[W�@vs�Q �v
W�����j¨&0t�}6�+��(�Z�t��}�8�k��q��W���-&�$����?ۜ���m�v�"k)���������D�1���Ҩ���#��7��=�G��|���d;���\K�l�7O,�W�Ӿg�X������pEd??��ɞ�Ej^~�a "�wD���oVt:Za����4�\||��My����gsDrl	$�t�ڢDSJ� ��sR��Ę�}���SȚ^O:5Ε�y�A	ݸP�_���b��yQԊ��V0ZW�I�@����E��DM:Rfz����o�i��L���֬ѱa�Z-@���G!���-���;�"!���t�u/�",��	r�L�����,_
a��?�������k�M}���ӯo����UT���>����)F/��hTR�֦�kH��d����y�i'0����Jb��mu@	h�]
[�BC�}zG*^�xTgb�$�~�Z���^�?·�L��C�߫�8<��B	_g&3(����u?5_�����IP��y��#F�͂�3(m�f���O���	�٘N�n�q�����(|�}���o��f��� -��~z}0�Dsf�Y�����5����E)y/LZ+_�N,2�[Z!k���j��7565 �䧽� aYH �ż��C�;��)����8�ře���6䇂���Ù]�.d�?����O�f��#�@'���J��=�پWo�_��z�@X�[57��l	
�>��)����~j��Q���i�(`s�8�E��yJ{=ϭή�ѧ�S�[j��;-z���t�i�@�OEpj%+�0��F ��!$�"��.�M��2�G�����8���p"��~- ���B�����zN�����ة�t-6%LdO��?��p��������z��Ym�V��\��_vN�=P: �L�,�T)���<Z��jM��9��22��bD+ޘi`�f���Z����^��Ra�P��8�,�ٚ,w(UM�Wt�ʺ�
���unf._��� %h˧z� ���Ǎ�h�;��)��������*�#2I�2��3��[����U�I~"@��)bce����d�v�5�O�Gx��](��KU
�_6,�@t�h�B�v�$7Z/C]d�a��?Qqg1r�Z�'�5���ت�z7�H������8���J���63у;���-�>{��'|a�C�TӆboŽ��3����������#��󳹅���5��_��q�1��2F�:� �Y)�h��P,�it�`��ح����uJ�k�+uW�P �㢺�w{
�������&d�`#L����#��P��?[H�=���^{�9�N�%ƣ��Oxi���Z�RZJ!*ԁF������ƌ� /g;䋯�Li���Q�5�{����OP���OA�lv�%�*�U�3���&6-WRa�c��Di��C~�}s�A9��C��:�MM�j��c�0� �D^r�� �8�W�8e��������|	w �� �3|
3��&�1�j��������z5��*�o��Ak�;)�i�=Q-}�M�X��S�����R�eCª�N��I�R���U�\������8#b�,T9��;1�-GK�
��=c��n0�/��~_�<f�P�aX�E`���Y
&�W���IB�; �oQ�Im)����"'�<����0���[�/�ZJ���3��b\ޫ��x8Pu��|@���ȟ���1���i�������~v�U���ʩ��T*����'�s�X��!!���q%�G��=c˫$�7����`���%K\X?�2�Gc���9@\s��2�z�,�)k�
Ѵ��B �:<�ӯ�� �L����%*i�����2n��E�T��� V��<>9#|���%e�,̹r܈e/~���Mh<'�;���{�c �fMd��j�$�K�|t&�9B�"vHâ��"�~8��.<��\���V��<$߇���,efa6Y�d���:����]���|�a��� ���r�t��V��oh{%ƗP@�͎	�mOPڬІ�,Ȱ��l���XuRʃtDJs��pQ�;���Eܜ��p*ٯab;|�UpI��
����,I
�ޞ0�ؒ#A���.aԚ��$�RĿ���@����1��.�� �aTa-��Hv0:j�Ź�W�""��V�\b�#KE{�J�2y����$�&�_K@���q���jϹ6-��`���ؕJ]�Ӧ=�B���op��9uAkz���p5�^�y1�uVgF3�/K?D��Iiєj�6�g&O�XFn�N�۳J����pc��ˊ�%U��%|(b��ҍ �M^�����( t�wxL�ߦwp�UUo��oUO��4:5]�H�|�i&Ѻ��*�������w���'/BSV�9�	E�
�F�8|t�U2� ?�r0��	�ѕ�"��1!QeӴ�0�^�~�F<i_���q،%Pӏ$�
����Β�	H������C�����Ι���ש��}��ꧺ�-�7���`Q\n\[��DD�@�m�l"0���؋[\j����%��GS`�W���m��i5M4��^�m��ߦ ˱���cW��o�H'��}�űT"����=
i�,��G�):�}�H�N6�N��|M%#�7e)X�*Ģ/�@���1$W&�N��n �08�{}�S�5Iʮ�sS.,I5��+�k��\"�
�a:�M!2�$��;S�v�+��BhkE���L��"N,�F?q�lx�;%�8���ٷv+B8ug*$v�+��$�"�Ԛ�V��Z�n��LԐ覸��u��kǣ'�A����{2�7��7���R7:q�w��Y���&Y�!)P�jc�O���R?�Ŝ��/�^K���{��<���C? ��r�}C�(������VĢ�j�Mz�3�X"�}�Xd�R��E8+��G��H�N�ފ�|�%2%X�?�!{�=vO֊#�J ��;�6_�]��Q��pݶ]+�1������i����� ��ր���@g@-,���~�8�b�n�6r���Wi��]��W��6/#@�X,%�Wp_����5�ܨ�v��C���ܵ��*�;��u!���䫳���i���P�&��m�LS����SYԹC�J�«�_$�{��sj�\����l�`SA�凖������Q�3�͗ϵ�õ]dd��7��3�G�n��oO�׈j�ޞaJ�jr�F�N	X�h��7�[��?�S��Z��O�>�T#��F`���O�S8�J���`9�-9+���bck�?iM��>Ӛ�n=}E����Z[�X��#�˔A�z�M]�E�p-�ʄ!E�ۗsM*�|��ʦ����[6��1c�ɢ@j��vE�X�S����X3����o-�� і[k�x�S2� =eS��Gz��HTd|.H��!�I�9���ъa���(];5��I�nݼ��~BG�C�jaG�����\�	�
����f�}��4hL~��@|ݤ*����Ӎ<�|p��7���P��D�V+5��{��n"6W��h��P���	,�u�>J�ճ��������rM���
MTU���n-�b>�m�Oã��I�gDn�Z�񮒼Ң�\ �,��+oz�1��|rX���L�T���3��'������M��,o�}�{W�\����x�L�t��ၿl?�=�Z�������d�T�]&W�۝���&
p�������*�l$����	�?������?�4�\c�y��/I=VZno�0�a���ҥ�0cR9���v�NS.���)�~+���F�ˑ!�?9���"��TY�Rӻ5$u����if��ZB��Xz�R45��jq�����t��^��Q����9b�&M��꼻No���3��=�Y$r��g�W]Bٵ�h���"�U�T��RE�UQ���1�~8�.m��sl�[�r�]_�L�ʃػ�ׁ]�/��nh����]ch���'��>Ns�/��ph��U�]��c������R��!2��\������#༫;_�/�@:^��J?��l/&٣>�v�T�0(Z�Q;��`(���Ye*pl�6�}#����+�C������1�j���d!T|kԅ_���T�K���/�-�2��{j������{:DӦ�_\M\�F(U�`��(ƀs6r>�j���]{�)���EsTsTH1oqw��{�շK *��zd[k��ϧ��]�>�Zڟ��K2T�rlڥYD�|:��_j�R��J=p�N?�!����,(�R���F���5�z�z�����f��&Da�KT�D��2ED5c_���	���wj��)����3B4�t8~�@��>�4@W[�O�)T6��]&�N|�B��8���n|^��5�8b	rF/߄�%������뙃X�t�F��Ko��d[�=K����nY!��������)���\�DLQ��&̿�9�&���U�-���	ا�]�g��H1��n���FI	u����z4I^˻r�l�$�{�g�p�/�[���!a��Qۮ��i�ip}�D\]�g�	#�2���������}����cU0��L����Hە*χ'�����)��u�K9�O��L�$8]�rm��[h@Ľ�Y��Y���2<�
<�gG��}c�Q�Y�YF�u?�W@��Y�����!�����ұލ�*%�[؄�,>��y{�R��ۍ ">����{�)�0X�?!��ڰ>i����cy7ug~���5��nXY����2����b%�{VIE������F�N�����gN�g���%V��x��8E"i�IL�t�WK��,�������؍F)|6��+Έn9~2�Ƥgd����=�ֹ"��~�p���߿a{Sr]�z�a"আ��Z9��L3ܛw�g�φ���(f\��-Ja�s�ʱ��Rp�+\a�v��y
9p�tP�,v���'�y�@̀SN�#�X���y� ���h�*	(D�B������m����iX��(	�V5w���2��o�,�@� ja,fj$��#}�r��=��R�_|{q����x�}�/,KL!:9�h��!�h��/��,��;8Up�B��gπ{ru���\_V򭋓@�pPM�:�az=���f0H�y��seG�cL�\
���Gc���3	~���]�l�����+\Ac������\�?�ff)M=-���� ���� ���֋C���U����	�-����7�ExDҘ~E�M��8@q`Lsi+ԑ��-;����K�wl��}�&��2��:q�G*����@ڜ���S�8&�k�Y>��f6��k+�*�z���Sk�%��RJ�	�P���D���usQ���4gW$pc���uڊ�KbUr� 9�%�r���0��Gn;L�rm�ڬ�:=�x�:U 
�|"E�Cڮ�fb\Y��;� �LW�d�qIή�P�D�$!���6r�U��+�:4���\���_����)���	b��֞�O�Rw$$��yw[�,%m�2����~%-��@�SфK��)e�#lb���D"_
��聗���N��� Wr!�E:S@��]��KK5�����m��V��n�Iѹ�~D��	�3B'q��lQ� ��ѱcU���D����5���=a����L�7~΁J�Z�> '$Pm �=D�����s�����p�7)uҍ����DDVz}�����%;X5���|������ȩ�u皓D��]��T桉�֑�`R�nVէ�V�����,��(]]�����(�O���|��/��5�X����5���F��_�������}�aM�16cꨥ��~ �$��|gm	's��L�tu�'�Q���;+"����ӧF����1Ac�@#a;�HC��PR����8�Ԫ�^��=�l�Q%�,*-���Go�b�����Pp�n��U�?b	�F����I�x��4Ӷ�;�p	q�&3xS��*bO���IX�ݹ���,z�j����<��~�Z�>l�)N�@{�Qބŋ`35�(_���YU����(�ޜ��A����[Ƣ�Q�{2�<��~��9V�d���k|���٢�8C���`&���9��+�����:�̮�$	�N.�\���5�hK>���+�xq`�r���z��w��?K�Qʑ� )��3��W���S̽,Nu �ap�ٗ����g�g�$I5@���i�v�|�{�˕9kD��]��i��\��l���h�@������2h��I�0��G���p�a~�8���Q*r�Î�|�#�y�v�e����R','d��Α�[�!S�x0��G�}��ld�c � ף	�o�h�f����}�[��:�Ȝ[)~
���~Pb7�J���x�A���X��S@RVr@���:=��3�L�+�����[*ĥ!@6>�W�����{z�A�n_�kwA}N�YLZ@�]���/<�O�Ir/��R/eM���N�&�� .��\���2~�P��Ϫ�I��Z��=Z�'�p����p�Ń�|Pda�pY�N���.������e�b�]����T�:УZ���M��h4J�p���?��������ɟ P��ٺ#>��Ռ���/�̧)]	+Z$un���aj�C����6���@���2e"3ׯZ�4[�(ļ#@��a��d�8H�z�O	O\�vo6v�� 7o{6�� ��:ʰ�n{���-ŕH����:�t��3��nK��N=p��3�D���./�`��-�1�#�G���ѱp?�Ȑ�\���Y�TR'�0���B�s<�7�@3���ˑ������ـ��t�0ظF���ԏH뤟2q^�r���]a>6g�+�m�BX�!M����[y[��'?���翖Nzi�S4h܁ƍ\C��v[��b�*��a�����G�C��0]�Hg2J�4|��b��	��;2��56iL"/?�+"Ƽ��%���G{�&<����J�2��Tv+��b�|$��e�/a�Ե��z-�2w��7f)tA��w�9�ȝꚓ� �x根�R yhTSΕ���x��2��q�Hz����4T�ə���������&�̀��}�^�U��C�÷�	�0��@��A��O��]!����*�p��z��㛰��ݺ1��|A��q�d;(�I���}t�4�h�(��t�u���B*،����z���AFuI��i��2_�'��hq�k��[_͈I�Ѳ�B�	�G��uzX�q�$žk�Q�3�^K�?�����J}�az�f�饰tt��j�^J�*G`�,�R�}H4�.�����S���h#�⁅J�?
�ZekD�pO��k0J����Z"e�9M�`N�2�yU�i����]H��� {�j�=��aO;���0�Dkp�#�¼7�%q�(�N�:��!�6 ���}7uR]�n�3�k.4�d�҇$
OȜ��T�:����Du._^V�0�U��u��adJ2ـ�s()�e�ip��3+�x�\�\�ep���{�GN5�������OpeI�Z������S���NJDZ���M���M�=i~1:�3�z��K�_o2C�t5�=�ړ8�4�u�%E� �'��F�� �^ܯ��Uz����\���h�#��������������9^�u!��fC�iW3ץ�#�.�y��z�բ��I��X!�������ߺ�6��	��i\�gK��{IJ{	��Iq��F�����Vq㢣�Z`��=�⤸�n��
3`;Eb�Jvc���ps�3�h"���3��R���q�~X��+���i�b�[�0���в���JA���H�������יߟy��ͷ�F��w%��%����(��6;3w]�h��C���~����y�庞
:N�� F�Uz�+C��è������H���`�2�@,k'�*ǡ�:��8	�d�4���|�(3�Ƅŋ;���w��I�$9������*}��d��cя��@�S�'��⤋ �i�ǐש�kl:�%b��m�oC�!b�d E�l��$u�_Ķ7�-����|i�(K'���`�X�R5E�Mk�i����lOЭX+�/�˛+�=���L�cT#�V�0&ĝ��R�-9�#�� N�N5���1c� �B�l%|N�֬j��Q��=��U�&u��S´����P�t��P%O߰�,\<��ܸU݄L��-2�u�ub�	�zl֖D�C�EX��}�8���/� �>��v�p}�lmJ!��]�Mb�����o �*�$���۩�3j]�O��)Z+��7�h�u�	mB�b褚�o3�/��H����I��V��|ڢ>\��5�z�"�w�_�%�mU�:[�2������{���
�L{?"2�>�'�p�$y�`V�?VSn�Ӡ3I�T��?��<����dO���$@����֬b�������QQ	@�E8s��UP1�R�S�ƍ߯��y��u��}���h�6�����H���H�HL���9�
��տQ�S�=o��M�{ڱ�&�[�/~I�h�0�Tǎ\��|�*q��`h�̱t@��<�7Q�xh%����ޕ4
Р�j�'���#\��l�D��jR%8Jj��(��^R!4`g���A#?#������E�3`�C,���M��	�(��~[brq^�j�>�2�����y'�׶ȋ��3�iu*��g�v���j*Ā��[<�Ra$�����)�(��9YF��'���3"��P�����Gъ����$��O~�kL�P��!Ɏ�6<$��ޚ@P���+Z�sl�<teφ�Q���S�	�L�d��}q�i�&�0�Q֡#�Zy�'2PP��^��+�>���%xh���Ү�,�+�ְ����e�Ϋ\@>`�RA1x�����PU�L��'j��q�IWl!9�ꅴ����cuj�niW�n����W8�c�zN��=�>�x����"ߵ��G�D�k���gӐ��i�.-�z���X��3gV��jo1��e0�~���-�6`�m���:�͙-�s�K5����sds@n�}�VΩ8Ԇ<�Eꪾb7���d�tP�P���YI�i%�Wh���<��}s>�o����r�U�0�0l˧� ���r�nu�CP����KYw��i�=�9R]s����.p�[�y�o�T��k�^�l�h"��	��n��5b6�O���\��������B0���ău���߅�7�i��~���Dx�+�N�L����n��Dd)����q�"Uh�e#�{��\�����toq�B1\��ׯ�~5́���Zw�<�����)����Zknw�p�Jq~]�g�;}�3��&{���Ս�&��R��wx���b��o��8��245���#4�D�w;�3n%������ؓ�$��/H(�&�-3����	11�LWD%�(��ҍ�����2��f��|���ڐ��HrQ��n+ �J%��(�J)Mz8�^��&N>���u���u�D0�)����f �I(N�=�dy��Ϋ�ZxA���p���F��-�����}�޾���:Аݏot.؟�9��� z=�l$����>:���V��w�����"�
����e2��|E �Nΰ06�@�7�H�a!	�������g��D��1��I��s�NYոY�O/0Ar�&���)]��Y�bl���6�}3�M�-X���\)b��h-l��悭ą)�5RoQ�FI���!Y"P�����s�{wU�z�vw �*�o�mǩ�C�8u+�$�r��땨)�+[2־�ˢa�J8�����ܱ�CJIgs�^�V[u� rO��O����g*�L���Ȁ�\��3���r���/�l�C�?���6�Y�4��8�8��Ʒ�3Uw�b4o��\�q)iEl �˝/��� ��H.J=���q%tI�c%E�*� n?�.�Ct��~�hYR��G�h O�*����<�{f�w�AQ'(�Y�z�oz/-�>��6�Si
Me�G������0�m�%1�V���+��]a�h��R̜q�V����*]���8�����Սf�bNf�a���`�����H �Vy���(g�xL�a?�:��=�t�����w�aW�0��G���j�7�d���x�{�f�"d^O!�w)��wt�O��+�4�_�f��j�Tk�{��� ��N��+՚���1�P9R�Ȕ!����PK:���)Ϟ�^棟���v:٘S`k_��)�����7ZJ�m	rPv� 6�i1U�T7B���H�Ϫ��|�E_ n���D�DL���`K�Z>��w�븮V�"ۣ�
ӻ���cߪ�Q�_R���6�_�Wkz�눸#�n�E���%��h<K���X�L�����cw	����V����$߱�Wc����7�eG��~�D]|�6� ���rw̒8/d��sb��hv�չE]�T�+�J��o�|uq��BT�1��ɎY����꾭+lQĭ1˧M����J�l��m�M�x�I�� ��|Wk��-�u#w�n&7��1B�lj��S���K �2������nj��q�;z��aR��Cx�N-Z?g�K�0��E3���u��1q���B-mӸC�U��è�%u����£p�,�Mm��]opMi� ��+�NpU߄ky�3��q&:%&�{u~f�~9��\3@I���K*�^�F��A{"ٶ/�I�p� �	���5����m�晓sc�T��	~ 40����R�H��0h�ɕ���"~�����`��#24!p���.�f|�D���'�D�m�,0�Cܣ%Z�8��"9H�q,�r���Ue]�f�y�*�v� �X�`֒�BA�py�yh�Mp~"0��������7lحM=��C��}YQZ���^;!��Z��-z?�K�f(��ޟv��d�$����g�' �r�qY�����<��
_�R�|�:�ޙ���Ư"~2�66F�p�lʪ++�z��K[D�w�l�
y�i�T�Q������q�ph�硲wޟ]�T!C>�q����]%9�NQ�L�O��5��HÂ|P:�_��f�FU�f6#(�w���]C���S�}	X�A���*<̽l�sJ½M8M.�ʺ�
��V���ʊȲU�Z���������g�
���@���/�Ikc�	Y-�P ��E�|���%MM(6㭥�.:H�7��Q%�rݲbT�2M�t�V���ǋ��u�/�_�sͻ�1��U[t6T$:}�t�D+���obz�$��i���}���`�����G'&������� �l�c��k�1��� S�U<d��ැj����#ϩ�9�q�i7�=��'�¦ov��i�c��	�݀��|�2�"*�G w ��|G�� <�����o����N_uƖ~p���\�A�V���L�Ǻ�-�vQ�H���}��T?��7��B)�ڇf�wD>j�^���!(zoL7��v`��_h�k?Gf0cBfCa`�h)p�D�k�~E�V���n�Dh���H�������[�-� ��r��bH����e������2S����^���*�`1��#,�o��(A�r�e���=ʎ<]��.��!��D��=l�N���>���wed�5]�*��eC����0�]�ݩih�^��Zy��X�i̬m�.ؠ���@�}�6�J�U&~�z��\s�10����4�no�Y#�]����	����$~����6y<f���s�x.z�Q�U{�"��VUpg�+'���Ƥ�p0�!�5��e���ɥ�_�Lq>��PAr�����*�y��,��	���nD}L�#%���g~f
#���Xꕇ�3���~�E��с�1�ЌeK�*�����N�3OK���ATe������by~+����3�9Ƨo��n��-��i��J�4��?�E-k|��_���l������m��X�M����f��-LJF�6�Vg������J�z���u�_@��b瞞�$ζ�a�Yr��c�g
�<����yv��I�(�}l�vLXW��h�-p�J�X'�1���&06�-�\D��u����@����jw���,�2�8B ɔԬ�S�������g�1$�w�y7���T��DI�4c�B����9� K��D)��:|
����_$}���mJ���3�+�O:�aL�	Y���������h��6���DD�5I��ӂ�T����s8���g�sJ;�����jA�J��q��e�����q3$��o�%�տ(S0���mBD'�:H���%M�z�īn)mZ�)f�wmHΆRuQ�/���/b�T�a#��l�7/_%�'�V���-+@�g�L�mz��J�]�QD޿=���'	/�i�S(�jQ5εe&8 ��Q3t�N���Ҍtu3
��;�tI]"<�t�z��m̽�g�>度�O�o�w!���8n���B87½&�����f+`�G&���1e��q:JV��ש3ڣ�t��?�A^�Z2AD4�^�B�٪�A��ҫ�Aw�[cW���Ц�XZ3�DH�Je�*��~�6z�fL���涼>��S��e���,�kj��T�A��HC�"��=��)~f����47�^0!@��i���ʬ��u�ac+�.ᵥ?�\3H��C�3�-�$�����~���K�o�!I��S�e����fx+�=+��M�O�$	T>MKI���S��~����<r)����|:�\r��P�ݎ/n�k'�e��#{CV:��Kt2�B!D��A���.���n�ל���D<�bn�jƢ���'�M$���x2{o��,�Y��$�)a����N���:u��ޞޝ�ꋤ�$�!��65�*R�糺a���eK�V,KZ��Dm��V��E)<�����R�4��'v�v��j��s�2#�y�*����Q�!���>.<�H���_�2��5��wY�Q֌��O�Γ:�fm���e�t$�T�0�{�7����
^�"X:t5)��SI��e5CBÂH�;9��B�"�������m��q�7A"<������X����0g��ޫ=��iI�oV���ҚUL*��i} GdO�3a�n᫿����Ar�e6�1WU��Q�n] ����KP��9��l%{�����	���=�#w �᧖�.YU	�B/���_���X��j4�KO����u�D1cu]�t������t�ZS����ĥ��R��+��הG:��!:F�h*"/J����#<��L}u�����~�S��#c�0�П��M ]V_�:��ӈ��	�ѥf>����;��ʫ5�����$AC%�'+&\��Q0 迧���V��� 5�n���)�"���z������;^���y��B�3�?��{�Fa�o�]=�m�g(D��#,���-��OƲS�q�.[B@��1z. {�o�{>�a\��I�$3�V��L�<���3u��,\���hy�U򽒰P=u�j�nB%��=�)���W>;���0#.a�*����U��7�r��޺2to*�+ql�s*p̦ ��ʏ|V%'|�'e����n>:� G;��?�Q�5g>��KTd��ǅwJ��[.Y@��ՠ�38�'�߀������W�����>����
gb̻�UГ6��9�s��o�����IWpTĭ����|�v�ۆsPO�܇do�öX�&nق���2�5��+ʂi�-8�n~iϲ6�2�z�� F���H�t//s�E L��,��`?J*�#�.r�d }J�T{��U����&��L�4�UR-Ш}Ӽh10�6탯K���A�Y)�r4��_*��Qs�3�G�x���*��1{��Rm � L�+��/����W��8��ȕG�}wD"W������l�V�O�Ok7�Wj ���JT����Po�U�^�~�<�J&�r�I���580�V�j�JPz���A��2���Y|:bQ/�g�$�Y]��8�|0+���� w��]��
|Q�v��Ai6��M%y��0�ìf��z����M�e����,m�CtQ���J[[r�7��3�O�1r
>Q��߾�	�5%�����Xw��� 5����jg�e�t"5��6�Z�έ��SB��;
65Ou���֎\.���k�mR������ln��C|����%u���֝9@쐩yj��4�G��ػ��o����������ѼfY�F�����5�Gгt����C*ģ���P�2C�����v�lǷw�>�n�ʋ@wy?�����N���&��ע�䝴<�~��]���;��B�^�� F_}��4��=޽r�.���LD���v���|n�h��Ѕ���F�����^p�e��6�&�JJ�$܌���ϱ�`bh3�I-=ު$�>�w���u>�~�)O�b���"�WR����[�5鳊�ēm@��װO&Ъ^����T���m6ÇaJ��`�4��>o���B����������L䃕��h��[���+c�w*-��ah�3�O=e�s6���U�%�Ո,b.�����c�<��Mq��S��"mI@��+�K���I���QW8I��
$A�'��7��J^����I����CU�Ԝ��+=���ީN:�Fv�m�?O������dLi"|��[��-z�3�P�3gE��	$��B�GR/!曣��I����1ܥ8�\��"�
0[嘛����x6wLs<��("�{׷�$�K�g�?��3���Tr��hÇ#ԌIo�1���͞kZ��zF��/\a�P�r��b���t;S�ń��M�t��� VE�>�S�w�ׅ����TxA����i9��~�F�!?T��ţ���U�xNf؍!���Di��5=�ɎF���`�uJKSI-���~����5 ��?g�l���M���*���hT1�!w"ƿ5A�E��xׅ '��+�v;��,���S����Bp�y]��	��lӑ�RH��r> ̮��[�9ԗP֒���,
H�˪Ҿ?a�c4D~8�f�~��<͔�.8ͱOq�x���d5���T� ���4�. ��%����Q�D�H�>~��]��j\�� �KT��2{gfi�1���I��Hխ�y@�p��Yf�]�6��P~Z-��{yQQ!�,~d�ŋjR�+@�s��Sh�����K�-F&���k�W}V9�D�7�E0}4O=ڮ�[�Fl�$��c���G���@��/��H�&��$��]{�S0�R�lH��b������;�('�����Y3�s��
�Ξ�a�Mh�&ӋiqQÂ{�IK������VE�J�����%�M��������������X���`������v�����^�ͺ��?g�.��>K�ǽ���u�f�B�ᔕ�3���T�JyZ�Ԃ����:n�b��H*
m荪+8����p��T�&��Q�C��oBAm�fD�}����q�[�6�!�֜f�&V�B��kR�T��ǟ�f�'ށ���.#�`/EfE���'�I��'��
zv�dC���d�Ob��jݎ6_$���Vg�<���I�8R $b����?ZR���eS�i��مN���� h�-����n���6����)ӳ�#�����k��?���nGFg9�>6P�+��Q�`�>J��nt��x�&��Ј
��=�2�אV^��8E����gO��6[�'��C	��h?�W%A#�%?;"�=äQ7dm�����s����Ɇ��G� �'�ҽ�?��0n��^�v�4b&=F��d������{� ��C����PǬ�X*�ټ�ׂq�GDw�{����E�،d�[n\o��Α�Ak���`I���ę��}���S�q7�}��q��.FYH��l�wS�Qq���W�4|���]��ph��&ž��R��̩2�]��nD k�����!M����:~�/��=���ҹ]�j����O1�L^j&�+��r�G��\�4B�r��y=����7�4�ya�&��l���!�}�>t������z�GaL�fX�}��J�1E�LV^`,Yu
�2�r@V�J��DGD��a@���Z���Ts�b�#4�v�����\��|��+LC�^j��f2��Lz���ƒ���j����B�Bs���OV݇�����?��a���q=X��d��K�HP��v�N�L�^/���oP�}���~=M�뇿ͼ�1�������r�3������� U��M����q�o���E�n�B+�y:�M.I�[�A��0�nMFSU	�Q5؟��]]Hr���L�p�~��WC�C	��e�ފ�~�B#~�mSg�mn$d�)$��Dr��{�����a�>zAK-O�1-���>V���ڋG[��hCBK��f9�*��2˙�%
8/�,���y���nD�m����;�\��H��d�:�w7��� ���<ĳ�O.�h��n�H�<�%R7z�L�n)��Ҹ1�2�a��|�r�i�y�{*4m��ة`�6h�nQ�#Ժ�̤�-` &E��^IUq6�^���4R��h9+�Ŝ	+��	o~<���H�y�.����I&����_�%��2W6;o\�m�q����e��sb�E��vN�!��Ǫw'쭞7�o�z�> ���h�%�sl�yqN����B_9g�����1L�Lo���u�.+�g`{Xetc����4[?��0�z��G����!�I��.nm�y����L��r��x�ռ�؜���N���ܻo��OA�ah����H`��Q�,��̻�MG�[�% ��y����d-&��!���gC���{��Ԛ�&��w�$"��H��C�x��G��Eϝ�r�sG~������$���M��Fǜ���%�Y���<�v��A*�v�:��1z@lV�ҕ.��9�&v^��+À��ݪ�?7#���X��q�nu`]Ou��oR��5fbA����s���:K�6��Gfẹ�̸�p�:~Yw�8��y��oY�`�����'+(B�x4��
&�!��m`��m�E��������9��d�9����0YQQ��E,~�xh5*����������#�"=�g�����C���=r�S���Z ��4:�T�W�M��k�O�n��z��h�в:�
Ɉ��a��X���<�zE��k,�?�6��m��aI�,s<�E]��Ϡr1P�?��*������?��^����.�,g�!�.vpi3�יo4)�$�LvI�.5J�_2"��	�3�,���Ⱥ��	-r�띊�U����J@*�!Cjc����$7ޑ���u�C�[5���1�Jm��lCV�?e0��0�vV��D�qL�!t	n�5a����u�DJ'K
��WпM����G
�)(} x;0U^�`��������-�
1�����X!G�rPG���$��x�q�{�X�@�eA���s��|���<�瞙A�Iv�����J�J5���M�{7,���`�򣜁o�A_ׯ��ܩ��k))�N�SoM;�H*]1ێQ�o�8�\�V_�kEx2\t�y��6U��|��ٓ��>��W<t���ʼ�",�F��zhq���;M�K��ynO��2_�U~����Z�����D[!hMj�B0N2����򋖛�I�H�x��Q���Ը�A���.|JbK�6���Pͺή�i�т#�N�' ��}��Rh�/���ԡ��P,���=��mJ/*��15u%;���rۂ��"��Y���-Z~P����0C��W|ez����{m v�^�ި�<+r2r'�~�ap�Rg"q�9�)ȑ�'�?M�}5֪��Ԟ��@���"�-��&ʲ���f)�؃�8��{k<�\1��B3�Aw�+ fyp���oo}Yg���4`��S�=<ߴ��!�Tg�-�㪪n�o�[B,F�p:�@4z�jw�uX���I�҄(��'U�2-���,�h:J�ևs[5��hf����ҚӸ٨����0�37�T�0�S�Yu4��9��6�x; ��F�������fs��<�|����=����l�\El��������`�����t�JҴ��W�I^���c�0�İ1��z���P�ن���铢��:#��s���~̰�f��u������7}Rg���6D��2O���:����<˟G��՜R�)��J3U8M!0왧��S9�@��'a޶͂b&�pXf� C�'Y6q�.����o��k2�$��N���
i�^��*r���&����4T8� � ��r�-hZRLI!mD��+�-'-�Y�W�4��4b��; <b��ӯ�0�0J�w����\6��e�H�F��i8>C����/lb���Rd�/�c�Br�pt�����T^���F�E}m꺦�X8�O�HLLOU�lgcP�%^���'�ݏ�3��Od`�������A�J魉̨A͐?�e�w��G�l�ЙǁE7<HH2�nӓ�Xz��ݭ��{��Y%���+�s�3��M�|a}���K�w^p��V�h��~��F��~9j�J_V��P��O���m����iB��ET� ՚�Mg\�b f!4�1!#r�C_�#��Lȵz��3�Jay�B�S�9!-!��p=��rOdx�B_YP�>�ԅW�K��AcX
�.D<�<\�S�gA�h�Bg�t���%&�h�51Tb>F���y�G���L��y����I~Q�mH��ێ6�i�����+�'m\Od�װ>��I�xb��%P���c�%3kQfT&��6-�1�~�<��D�҄J�IȬtg=���w�x��#��5�K�w�d�^7���;�`���z��0�TM��f�Bo,`�,�N�\?��
a���[�!�	�=���Dl4�\���v��Ph�����9֬@�D�b4�~9��UQ�j�&��ɡ�w7�i_eH��z��6Ӝ��>@����5�]K�yԙt'\/d�0<�=bs8��>du�����W'�yD����T��iW���|����R��/�9�LZ'�L�yJ}X��\N�+"�;��܆� ��
�O�n͵]�w<Y�J��Gt=��㟏j�[0�+ot��T,L�˙�%���>{�]V��d��9��6�\bv-��Ytn?�h'�4���hKR��1A-�*�&[��D�~t $z79h|�a4�Y�����_UiJ�Ӆ!�YQs�箎�a��WNj�^d�(DS�y�z�j��Q�:��ė:��C��j#�aE�G�b=�kl-芬 Ro6��]���z�0)����~?� C����\l� �j��#o^jS'a	�!�uY�q�Wc��7Ij�ٝ(�&�(t��-�F���)�?�ά����݄.%9��	m}`?�O+��yY�eҧ;N�v�B�IG�{N���L^���y����7~���a(�}��yu1���*�����ײ�1QN6<QD�j.3���V��!��r�X>W@�ݠ55�{}��f���?wN$�q:��ًƆ~��{į����^�0�O�ꋉ�n4woq���u��_�k�K�:�Ĩ��S%*���u4X%��L�vVn^�5Z_�5�3y��A�t�ClR�°O�ِ��� ".��d�Ԯ�s�� ��=]���8�^��s-�Eo�'~���1"郳�˘�}H��\�Ɉ�O����z�ri