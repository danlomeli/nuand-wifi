��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� rā�SZ )����C.��&0C]�-��[�3�-���+��պݣ�k�J�vo`�A�����f����u�X���v�=�а���]Q�Wۿ�߸�=_Q�X����j>��Zw�K��SvX��ƥ.���#�����Z�0���#7{��\S$��@1I�QX~TQ�E��db����۰� ���>0�%�9�j汈��}��1� ��2���h�G��SeY�a���	'<x�p��k�H`�H�j^y�0�s�78+���ֳ�`�R3dW��_��{p[�?$�s0��#�zS�_��bH
�c�p�IL7]� |����Q�� ��Rr���=��E즕2%�����`�^��l�q-�]�p��jf��Ӽ-f%H���ȳ�>��+���M�71��4_�) 3�46h�rb�J�W� k�h~K0�>P$�_n)���5�r�j��W�J&޴o��$>��6��ŀ�;A~<6P��K�~��f��*I
�Z��}`q���ApC��n���g���3��-�іrO�mF���,�$��@�BI�q�}��Ȥ֐����î�䂧��@������U���vU������ �T#K@f�㯁����|95<@���+�-�)�����K���FI�k���*@�m&���
���ma1[�2�u�I�\�U�yu���o�|��2����;�W�W�}P�K>%5�'�8���׫=����k��,�t�M�0�8]q3���N���GvZ�#z�HM���f5�����;�q��Pj����H�L�}��T7���z@�o	%�PFmy�lc�
)�8yIf�o���Z�"4��r���o�6˦��)��"�~���6��}�pY���]��
��K,�	���1D�̹�@��$���(_kk<| &���x,�u��Sm��Fģ	U��U9�k-��c�KU ��1$k�):h�����!�Έ>�l�B2A�V쉀�#� o�Aڐu�Q�%`��ܸ��cb.�����E��&�Ѯbz-V*�E���bnjۜb>W���z�<\UlA"���i��J��Xj݊���	p��k��1O:�$w%�C�\��H��U���Z�W��k�B�E��d��/���|�0�=o�g����/Z^����X@�N �Y*E�M��j��Ʒ�G��V��$��Qhw-J���,�B�����>�n�N9+���̍�)ТP��yw�~2�]�4�E�,��$&�_�������%�#P� M����PA��[�Z]�ϒ=!�ܠ��T�X�`2s��gq�D���&��%�?�Gy���4E��[4�͹��*�r�S�Q�����!P<�g����j�m2W|���i�:�?���_7��[�@k��v��I�������,��u�T�䷏Cë(��5<-�����8J���R�[{{l�Ijt�d�	0�:�K���}�� ��@W���D���&�b�kݿQ<
�d�dl�\aJ�n��En�V���pT���u!=��$�Z�
���Ѭ�!���w�*� ���NثE�_ *X��F�A
^�7��u ��*r�ܜK	���7�,+�iպ��z��<�7��x�j�ԡ��ܿ�bx2w-�lvDd�T���$:�k��l��Mr �n诗�Tcpb������/��h&�=��|�B"����Yb�=���t-�B��[K߹�zKVX�ʳ���_N��hF�Z�3 �<�8�=�yN��
��29b-v��i��4~����o���3Z��9�ӏ>ML7�"@c��"�nF*YC����e�]TZ����Z� ���7v�g�H1�".������	��L+3��J�a�_ɻN� �л�2Pf@OW:夸WvˌT�g�+2V'6�a�B�L~����@ƧƤ.`c�Z�nO��M:����k1)_����ě��`}��eU��	��O-&*�6�Í��.(���G���h����5κ�^T��s����p���y�[����nJ�c.:|]P��[��К�%M��h�O?�a8��R�w-�g��\j[���A|����a�ؾd*C���#�V�g����;��{�djB("��o�.�ur~��9"�|N�P��C��(�Ńz;[���Nq	��5S[���2ҧ�p�EL*��Op^���!����;;?�D�lJ9�h^�meF䗎[��'�9���=&��x� 9�!Wb���Da(�%�N��L{*���[�P�"������a7�e�mʶ@���7�K>	��B��Bm�d�̈��.�$)�$��gn�<j�}aF�μ���D��3�@1m�k��V�Y.'1�� *?	8�(-�6�$�/;d��̟�����5� �J����0��5r<��J���b���Ke�2ЇDlm����#Y��l�'����L�,�!fS���;���e�
�[�>)D{cK<p.����j��a��!���i��?�����bPr���������xD�B@Z�
Kb	��Y��8�6���,�Khc��F}W~x �����Ն��6z�����4z=�a�§��`���ǣt%H��@��D�pLQ���);��pM�_`}{ѩ�J5{�Y)MP*`�W�䚳?b����pB�DC9؇��_�sC����m'��K;�n���X41���O<��[Q4��ÂNh��TG��P��乭��iq�,�|N�)���-�<н�G����ܛ�/�z�E��,8�@�5�����e�BkW��)��+MOk��Dhyb&ry����r�C<aA�v�e+��t:?���$gr[���Ey��`��h�IW�G).��Z�+j {�"3��\&�����^��w�7�%��nҼ��+C��O�
'�H���ٯ��L9}�g>Ҿ�׸'_��3/�b��j�VW�%e�,i�7U�cR�3%/0��9�jy�S��q�b�*'"���æ���˾��3�%`��O��^��S6��$�5�tz�M���ѹ���� zB|K��i����mX���`Ί��iZ*��+�G*@�E速��%�<a��2:��n��<��Uk��@Jf�*�d&U|N`���X��n-�1����]���[�����˿��}�+o�R��	� �RX�����jkNaXRTI��諸*4�z�)���\�|?4￟&�t{��҅���*��>��3.-���rw����bV���I�]�aCF�dI�P��$,��B��"��d́������L5a	,�I�J�1��&EC���<�"�UB�Vy��t�)]�ݏ(V;��7��KO^�5�!$�H>K;E�����OW%�/��NÎN��p��;��5@u-m�=���ٜ�f�U��#��f�����>f�dF�Te�,��R�"]�۞U����.�?��*�!���{˹�I��g	a�n�~�9R�k�߂ ��(]����8���@��Jc��3�,�I��� &���Q�#w�Jv���K�٧�p��h��U� q4�5�^�*,j��{$���r��ŎD9���?������Ɣ/p��r&-WBR�IZ�E���/�j� 5)D� �oS����F��͛Ϻ �<s����f��R��*��_���<�38jc`8Q�L����#�_���W�6�qU�mX�����ƙ�lI���K=<�Z��|���oc�`u�����8��&�?��|00��H�{�����Ͳ��������;a��� ;��T ������^��李��rfd�0���p�.9��[�\/�A��r�T@lp>���.M�k��C/mV�:+�L�F���8�{�A.0FmaB�ʮ*HO���0W|W�x[J���P�f
{���o9�/��w
��ֺ�G�`zW/P��(��-�,�3�1H����;�?p��Aً�Ȓ���x�˿I��Vb
m����+FxE� /�a�Kt
�"÷��f}�T� ?^!f��d\��5>'��;��+�<�mt�)��,�V c��=�#s!״��\?)G��d?��z�랃1��nFү�9���Uk�9�5���Y��)���l�N�M���