��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� rā�SZ )����C.��&0C]�-��[�3�-���+��պݣ�k�J�vo`�A�����f����u�X���v�=�а���]Q�Wۿ�߸�=_Q�X����j>��Zw�K��SvX��ƥ.���#�����Z�0���#7{��\S$��@1I�QX~TQ�E��db����۰� ���>0�%�9�j汈��}��1� ��2���h�G��SeY�a���	'<x�p��k�H`�H�j^y�0�s�78+���ֳ�`�R3dW��_��{p[�?$�s0��#�zS�_��bH
�c�p�IL7]� |����Q�� ��Rr���=��E즕2%�����`�^��l�q-�]�p��jf��Ӽ-f%H���ȳ�>��+���M�71��4_�) 3�46h�rb�J�W� k�h~K0�>P$�_n)���5�r�j��W�J&޴o��$>��6��ŀ�;A~<6P��K�~��f��*I
�Z��}`q���ApC��n���g���3��-�іrO�mF���,�$��@�BI�q�}��Ȥ֐����î�䂧��@������U���vU������ �T#K@f�㯁����|95<@���+�-�)�����K���FI�k���*@�m&���
���ma1[�2�u�I�\�U�yu���o�|��2����;�W�W�}P�K>%5�'�8���׫=����k��,�t�M�0�8]q3���N���GvZ�i�+ C�e
��Ќ�S�v<%���q��e_��
�k�夞��>ZO7E~��5k�TW Aod��eE���G���ɑ-'���?�G$����ќ����8ɸ+ 5ʗ���l�d��,�J�
�^�3b,�����J����#n�zK����z�&��;|�\�^���'e�W�����">�w*	FO�Δ��v���I�h���/�*n
����N_����\͓O'������U���$�������es�"�<��)S#�}��o��%�:�mk�x���&�&@O�n�������cBT�Cb�	c+ʑL-�Of7Ug����:����'bX�0P��o�N���;6f���WѢ�ṬIB�&}��q��~���X�,����:�t��ߒ*��
��X;9c�1&�ٌ�yb�ev�bGMj"}	��ԛ Yq}�ￚ��=Z��(�i<u�D\�ʇ��1��,/�"UiZ��_�:T�9YG�r������+Z�N��C.!��1&�̲�@K�5�6��b/���,��,��--�ؽ�j8��+�kϗl�;�K�ޣ-%i-�2Y+%�1���ɻ��.�2�{���^�1~|��/Z�&wF�/%2qly]b�Ы������^[Ʀ��Җ�.:'�K��e�{�{�Eؚ��G����F(]�SEW#'{�z�̗P���������"Ea!��O;�V�Yu㵱�v����5�2H����x&��h*֋:yǛ�0�����hI�m"�4Y{ٗ���L(�+D�ur}^!
�}2����p�\�$����A�rZ��>7��������jP�z_����\�E>e})��w��W��ƚ�*��r�>b�wr8�V)v ��Ff"�ګ��W��P]yjc���&�o�`�U�7%�S@�&��W��ʊ|��jV�W.u�ID��M�Y�'�R䧣����z�;���E����%5�Z�US��ޗ� !e�G�!Y��_�'u@/<� ����A�D&�� �M\�%�aZ�m%��쬞W�g�jg��S9F��7�*����y�`4����q ��� ��}�\I9^%��E��z�ȧ�"�����}�Ԯ�G��8�k��=��\]��u#�+ #	�A�T>�ɇ�@hc���* �(�Nqyj���9o{��������1�P��ĤG܄)�W�Ś��y�|a���<ێ��߆�\f�8}J^�2hza�6����M�$��Ǉ���_.���..��I� &�H5����`֞䔌��.��lo��E�gpG���-�⺁�����P��6G˶5�UØs��	 ($L��y�{��jAy~}]�LA4��K�IA���6˭�b:�����y��܃f��� Jh��NWw/����@�6{�RY�[#%#;��O��O+U��q��P�z$_�Cѣ0GSP���	5��)�@8�}�����lӹ�����Cgb�u�$^�p!��:*�i��.�x���W6,�K�EP���Yܴ��AJM���6q��h�\ӔF���,��+(4IE6t�>��HN���x�t xWQH `�Ê>k�?jޮƠ&��g������[��c�\��b��h1׉�jk��c�	��0�?�ؽ��y�i$Pl��9�
�>��ċF7��V��S�U��J�ʛj�n�I�O���a��\��\�=}	���̧��O�T3ӻ���#B�{�E�E��`����}�SW,�\m}��eg�����Ѐ�<��g�=���LJ�;�]�� �>Dq(��9Ůd{������QP�c�]����1�����?S�y�$���[��N���?l���EvxϘg��&��4��v5���k��x-�ꂐ\�5mo��u��;_���1�
$����8˞�O|e�I�XVi���w����ٕ׈��_2��|��*�[����K��++1=��M�F��$84W���+�<�q�xD����#3+��Wz�-i�UO��"����p�2��e�I �����*h!ªl,�&���F�ĩ���[dci)箷LxҾop�znY��)s���cZ��Qh�g��J�2�g_�P�mI�WQ�mV`
�H��N��ft-9��e�'�(����I��jZ[I%bn�C�r�U.�se��O���AY���ba���#c�djh��M �T��Y�*��8�0�'Gw�3���4��q2�b/�Z�F5���ѝ�΂���$Z0�,B�v����<u�aT��,��hF=��Z)��8S�Y�5?X�TX�T�U��ȫ��ǝb{�ϥ�<�S�o�$�� ��ĥI)
���Ʌ�):����E�����U4�pHjEN��U9[^�n���2�-2A�Y(�JkY����_��ǉPz����9)`|�r
�8A��wg���Ɛ����v�E�ZG�f�V�zF&�P�64un]։��}��Ӆ�lq�5��}���6��w�i��93�e^C��W�U�ܩD"�-qd-�?���Φw��X��敖��p����*�� �&&=g�=v��E``��VC'�S�:����g�}�k�����.��"	�&���v�9��̄]9w2����ԃho��,��b��66s�����|��m��u����)����X&K3^b�Pb̵u�:�I#ڱ{�4(@�$�tK�~d���O���n\Ѽ�EPOq�f���PߜRCb^�s�=�м�X����3���ڧQqK)6�!��8!/�h��0�
��K��Az̃�pv}W� �^O���4��ϞҼ��L�k����w2�a�Q5��Ex�`��O<I>���ܧ<G��*�{J ��
��IM��?�����79f!jԇ?9��� ��~ĶxX�b:��;�Ѣq��u�Uc6c��ɮc��\m�K2?BL��L��UW���(o� �I���:OL���V4`�1T�}5�u���s[xK���ο������:�dG���t��lr���T�ʺ	�l`	��"�MG��i��I+��4���B�#Ar����:���q�}�= ��!)yZEI��;`� }U�m_N[��~(�����?�$>�5��sN㟣1MQi��]�%O?�2|����|v
�khy��'�"�`�����D$X)����`�HW���{�wY�!��%&	^��$���W�*l��Q1��=~�38�P`^�	���sS��<��z�CQ ף��M�S�c��r�� ׅu) ��40�4�Ķ��p�������K�e���(�ۤ�J��������ʾ����cz��TP�B`X��&�v��������/+��j�ڂ�=����?�^�2�m�����]+c]U���ڪ���J@���՞;ׯ<��!�ν}9�S�ۏ�+�v�(U娩���yךt�^���UW��85�1�������f<��`��t`��PL�Q-�ɼm���NEbz!1d�gb[�?�X]��4own.�q��ؘ�ٮ}Ӽ�%4!�pT��׻��vf����[�}~����s�0/΁�^OI#�f7
NB�d|�~�P�TϒП�1?Ą�����%���>>�k��.,7t�Vy���)M|!�����1vuݖ�~�X��4�T�ښ|�eD��_ע��,�v"�m���^̈́�����77o��)�E%�p�	$;���r��x��gq�%b���@�cG������Hv x4j١fD��ts���S�'-*�Z:�G;q�F�P�������� ѯ5Ai.,UE����B��r�+ȤB�^�W�E�U; �m�넖�(��vb攙H�F(7����"�N����G���{9HЇtBhjG�����]��Ǳ&��H]�`���u��ȂW&��81я�2��=d��0�@�K�
�~Je?�Q�ڏ1S�N��Pd!z�'�?M��<Up`���̿�9yK*�Ĭ�	"�Wػ�bS6��~�}'�H	HVnK1��u�����liD�;w*2��b��I��K��9t@o�������6t�������d�x����s5cz�rp�к%MuRY�QԸ�(�d�F��~&�H�xV4V�jW���8?�Ss���t�ea��ܜ�V��>&��`�.=��`�fg5�MjL���3�+Z��K�)'33�n�u:��6�͐�������f���C�ɞ��Z`���-N	�K
)��cdL��;�[����Ka���Qp(�FWMq
��9��П��HO�{!���8��G\��1�C|����` a��G�6�H��1��5����ω�c�6��w��D�=Z�=?7l�N�-]���$�'�Lp�C2�~�&.������P�� U�����ǵr��B
�)�k��NB�X��.��Q�R7��'pod>���浒��=sakj��6���p����"�d����g���!����Mq�]�'�,l����<� "�72�ͥB�M��p^�>#�x'���+���������/ډ3��0G^|��b�H���\������w�፨>�[ӗh��թ�:�p���^S�4�jpy�g��R&��[����@�D9���&��u�I
"�3jD	� e�2�*E*�>���R��m��{�P>'$�G2�21�]�/���J��Thڲ��;S�\��X;�TI�7���B��{�*&D�߉�-����T�4`Gau�P��*6=H	'O#�マ+_VA��:ƤN�x�y�����w?+-49����'�VK�������>@��ן<�[T2�w�
Ky�("��1ߑ�R���̷�"���O�ݯ�`������'�Q�<yjq��^S�-h{�9��d�4�]iS�)�*��:mI�CVW*gFR7
��*������墚�z.)�3a����fd��h���	�%|�؟6�Ń��Ɯ�vpٹ�0�X�~+� hGM�~)c����=�Y/w�l�N�n����w�mr�70zº��I�7m���ii=�ܪ� !(-�m3����\�!�N�y �X�d���`�ϓ�b�J<�v`Wʑv���b��b�!�x}l(0R�j벢�L�p!?�@�����A@����W��6��=*eY����}���6_���$Z㲩O�
q��e�:�VrlwT�\pC]9�`&��z�"��x8��j��QNL�O?�R���z��/���gB��%�kɏ6t�'6��Cs��ӝ�}񜜈1H_ޮx��h�s��$`���1/:���^��d���zٛ%�_��!w^㡹e�僣x���B�N���7�b�R����t�Q�پ����itR�ST=��爪rL�G�E����pi�`�J����3�3�0�g������k�4�O�`d=pV��;�>5:) �>�u���jU���s;`)�;����piQzSw���C�!�l���y�L�4��Lܰ�ƮMV-s�\�zpj$��g�W�25Ь���4�Uю/
��T���u�*NF�-����S����g�����-���B�dw�M���ђN����H�b����+�EZ�@9ۍp����.]+1/\T�rX��߀���L����"����� ����P�2�%��kD�C�<�O�jƫ�!"w�(����������֡���j�A��[^3f���G�O�r��G2�����J�o�2|$h���lKh��5vp!(n�o`jф�:�4C�X��;��L�v�O��3S����d*l���9���{�^�������¥�osO�,�f�k�6]'���xK#[J�0�<U3�u)&HD#�-=تN|	F�B���1��D?����5�.mPN��@��f$�T���R�V��nK���p���n���|���<�UM�LOGk"�N�ܫ�����zܣ�8�;f��l���a��\1����/��
hoa�a��M'&�h���������y"b�Ug��CGE��6G1K\v%ʬ�} %��т��Q�Qn�l��z*��i�]���g��#�[��7��(�|��䄩v�<�Em�I��/��<i�x� ���O������kD����L��q3u;$���%W�C�A��Ge!�%ͻm�n�M�&/��dW8�T���Kg��/b B��%��v�L���$��7���O�$\OfO����D!+� ++�a��{�:�&��NE8�Keý�NY���*J�W�4'�;,ʴ!%Tg|��c Ðro�R���4�1�3!��㬋�$������.���#$%���Q�M�O<k����Mp�i��@����e��} >��~�#yJ�L��������Z�J��	�jl��'_M�����Ѐ�s� WЋ��-���;���4��ci*,R2�I���ܾARs��K�fz2�_!fQX`_��0���
�I%f�Gl*?�Ḷ���u�.7t��c�$�k��G�p�z��e#1��̇��s����x(�;�"�J�ڳ�hf:��OEV��
�,n��C�k7���o����m�|+�B ��5�����\<O���O�M��ﳬiԙ�{��w���+�Ӭ�5݆C,��v*]������z�C�҂�U\��b�fv0o����9�*A�߼��jM��:0
Y(Մ�r�~SGZ��s����C�@ir��OF��`S�_��(z���O�g���/
'��ښ� I��[�d�sv�3-���/���Y���`^��ڌ6���M�����\�E�$�A��,t�Bwq�ﱗ�ω�g�T�=f�Z���gdLrŵ�߭����$����6Џ��x��ny��}f�7��=Ey ,��[)��e~��]E�z�R51Ƣ�rR(�V�M"!VÿAݡ d"f��jG&����89����r,Xy\e@�4>r��v D�˲����F�����-FFT��O���F-�-&���8��l$3�[�0�O? � �����QPn��V�~Y�����Q��J�i�b�,e,.�+�j;o���#l���eB�`_�
��B��*�)��e}qf�k�+�x |��`�a�$s�����4��Kx�8��Qj(2���on)��筇30��P�TxxV�M�q���n���L&�;���lO�֏׮��x��w�*8�p�j�}R&�7Ep����p,��K^��$�� ]|>�f��Q�
�����߰�@�8�y�Q�I�೿u�Ŧc-�a�՗W���q��)��p��L�V5�S�˳p�=�F��t��}�X�9&P�9$a~��=�]�H��
:yrc�1����n�j�ZXpy�"V_���{�eS��Ȥ�����&\˘�.օ$ixg�����ꐮ��ݕ�����p&�Zd�>|=��F��h����Aa�J�*����Ƭ+�z��_�^�b[�Eax�Z��8�߱Z����у���0 ��N�BfF�� C
F.?��1�JFHEZO�㉫�&��n�w�CѫS�sK�LX�E	�R��tC�
5Z��B�Ӱ�� ��Sc�,YY�UD2��N䞨s�����%�jƺ��gG^���:%����HnR>����8�H��(F2(�������ɸ��,�t�������s-�a5�'��ex�!*�$�j+�nr�s?��
ߢ��'��I�g�#:RO��C:���s�~���.�'�h���ҙ?��'���¶\�N��g{�F�/w��TdNe��e�b�G�ʗ��3gL+�u5�]�X�*�U��T���h2-�IF�+%r)�����.�]�"��(w
`!����rR���|���'�J91��3��cfN�/��x[v�p:�A,���K��C�'y�熡�R+�t��-.�9��t�����σG�S�{xZ����i���#9�~�ʹ��&�+j��j;�6}��Wsu��OF��	\��ܦ1�	���5,3����2؛�~���)�8:�u���c�PL�uQ�Zy���Gy�[NW��W�0ba�Z#S���*2����$�*��������`'�Fj�3a^x%Z�,G��ā�l|6�z,@�O���?�Eӌm��0M�T
����H������4J�ʱ�c+er���JbB�?���b����$�N�)�	Ōq,g����X�F�T���'iD#Bp1�b��h��� ��{_s���Z('lmQ1�O�ǵ�w�;F���ab�;� ׏�f�:(�Xu�P���ʡ�Y@Ñ]�.���X���ַ9�s�+ �=}�_n[��)˃��]e�kP�T�x,j��a(
!��g���顊���&�.�v��P�b�Sd�L^󉪨J�pT ��]'�P�FV�'hcp�Ї9X�Pߩ�=QO?���Q�锔~�	���V/L��Ϋ����0N*��L�.�H�� �A7p=����(/|$
1P6(���̎e�1X��%�����La{��X���E�؝V���AL,����lRܖ�����r3�Z:��R�JO�y� �J����7DdG[��|�?ɹ\̡�_�� ��A3��J��M�ԑ���-�|=��\V�2�W�2x�m6wX�)��_���9'r�g;��V5lYc.�ԑ-�!xWNx?��G��D���I�6s L��;���b��[�Y ӭP�N �ݪ��EF|;�l�j��vOb�Ċ��������Y��6�Q��V.ڗ$��A��_oJ�YvzD�p�C�5N&U��؄Jf�S����Y�X�g�~fm�V�9�s�6۴�徆3塂d�<%7FU�~���A�
>(�5�&���'B�y���FA�0w�m��S*�Ln��i�ز8��.��~����Z�I�yd�t�P�:�>����3�`i��ۉ_Zu=�|���Ba���b�`�kA7(U�'+y#s/�1�q��B�o�_�����]���=[��)��o}���"$�Q2Q�RN%���Y~*MPh�<��k���'�@�_�Gi6�e��0V�@3z܌�Es�}�D��ߚb)�Z�::�[�7�iQuq����0Ȭ�bA�Gi����+G�#�?3��X��an��QW4&G
�#��>����^����Z��K	q�i�WU���
0'���X��1#�D������`2<�k�E2配&j�TC>ωI{ k�bAdi��t��t�4�SӋ���{}���D�\z@
O.m]��O�Ok9���	ܿL&��/�9�H�R����J�[���PU.3���^Y+M\�!a<ުܚ�3b+�>Ƹّ~^�1/� L2h���N�e�NL Q����.��pϚ���+
C\L�������@��uJ,�����d8}c�iP��я�Z�������-����,6*��;c��Mb�:�q�o�EoA㞄�|��1�"MM,J�2BK{T ���W6�M�6��B���M�o�~]� t|R�a��G��q�\1Y�X���/��_�C�A�=x~���N���c|��"	JIk�=��<��K=�z5tp�F���Ss�GؙI��lJ��khZȣ��t���4j��B�Xb�eg!؟MB$��~��L5i��"Z�`8A���*��6x�B�9�u'���=o�?K�zN~�mi����u	�9�	�۟$`�J���;��2T����XlM�l=wG�=�
�h�x�j7t6C���F%�q�) �+��+�4tj0e
o�б�P�E�7_�N01?�<X�@ףF�qz��f|fڇ]hq}E���e��I3��~��r���k���|B,xi��B�$/cU�$�����E�y�d2n�+��q����l���%�٦0����)x#R(]� $7�V�H�5��x�}����1[��,i]Y��V-h��ke��~X�2C�zv��A�$��8H����Rp"�.�$��Z�²qL��P-�):�H�sTo-Ll��D��|���(���Ȫ�p4�+�*?&���4�&��X����<����]��SR�*8��`WMI�-�@2�V�C\H�h�iK���v$�Z���R����n#��]*�@m�)�h?"��d���MW�����v��ͥ�P���/����=k
��{C�P���^5���r-dp�K�ݗ�)D�1���#��P�)t]ٵe
����P-�z<�4L���ǉ ��y���9~l�A� ��S$E�"U |�Ӯ��g���'fqǀT��M�ԞIŃ�Zpʑ+�W�T��+��;r�dl����m��~GZ�o�%4Q%Ko�Y>��O#Z�l�]Du�Rxä�mSX�k~g�C��h��"����S��]��|5�c�-�5��ԁVvN�-lL���8%��[�Yj�r��1�5�j�d�WgL�i+x0��� ���)W;h�`�7@d�Nt-t�a�ҮDJ���VI��ΞR/g�u:�ak���ж��ì<�z�D��k��x;;d٬�]q�snY|�g�}='S�״v�?���`:e�6$j0(LV��<t����*$��sw��������*5k��X8����ȷ[_t�8��� ͷGA	�śF;l���D굳�y���D��B��¡�f�����2��Fb��4d��jI�r�����$��>+WQ�����y~1����Djϸ/�jLQ"�e1���91ʘ���?����]�#�Fn^�P�<; 	H�o�:2��i�V�C��-���;�?�����j�#
�ҝ�\��N���{�e x/bñjm9��s����ɺN�B�Iެ)��V���;`��Y�����.�0gŮ�2f���A����/�r�y��� &u��T�6�_'��޻u�m��S�Ӳi�
8>`ϋ�9�a`rǾ`�fZ��YY="��K9��43xjb�������:���G�&���y�N���HcO{���N��ȭ�"`�����*[�t�����@�[L�'���i� %i��7��s�K��I�/A��0��M~���2�N�c� G�5*�x'�Ō[ac��K�s4;��
�N���CL�����P���`���B0e��%֕��Ʒ�JƢ;�G�!)�&�e�h���V�Ur�k�L#ӎZ�J�Cy�}��ZD����ϻ�A��$�}��v����'gSr��+q��9d�3@���az�������Zp�ظr(�VvD��uQ���k�����H�o]�'�8�?.���|?ƨL��qk�V�q�|��������"h��:�q[X���0��v5�p|kv"Z Gҷ��;����䈉*�t������[��~���̹����饎$ (�^��k��n��,z p�f �m̺��冮4�g�<ϠM�o�"?8P.]�3�Wю�~�"�_k�Q��N_�q���������S���g�����W{F�O��eVT5n��.��z֯���(�Af^�4�-bGP�g��� ���G�r�b�N2B��;��d�q�n�v��?!+���d%f��J��E64)�vU��z���n��1�f�����5t,�,��M� 2��q�WܓR0B�\���po��;��_��O���(l$�,�9�`�=�w|�;����X1bx6��|� �ܲ�
"�R��֬pW��@��m��w՟��W�6�P��,�P@{)rы���:h���۴� ��E1RX�!/�ٿ�#L�N��+�)(�����dt IF� u�̏�d2h�~�TH�'Dϯ)C����q�����M���lʆ�yZ�jB��4�7�Bg���ʦ_g:������z����
3��G�W�ԃ�-��{�&q���+V+&�֝>��f6���`�^&��t�ۇ�e�x#�\F�/܍/縤���
?/��\B�m :�.
l�h`��	���x��'�k��m�^/���G<�>����R��ß~1����j�,��Lz�vd����=����������J�n2�U��S�]�!�������ژ��J�ٌZ}�6&8��~]���1�)���D��0�i��$N�/�O�(׀YȐt�KD��/����v�Oc�3Z$R�W��2�YNj?$3 Uk�\��f8-�f���;�ZZ��tj�ka1K>�D¦x�k������@�IKB��E1s���<\�<�p-��<#FUU0���/u����33b}���&6�B}����$���\Tl ���Y���ĭZ� �@���o��5�����5�I�go����]0;5�}��s#�Q��}a��G����g�`���ˈ��gF-�Q2.G^l����UfJ�).R/s�	E,�W�4Sc������I����E�J*�@'q�(1c�XV����%����e?F[A�8��G`)şq4]^�U�VRɲJ[Xd�K��y���[��_�0���*�,_��H���l
z;��4̽�}��4�'�����kM09�����S�=;V���=Y�.=�U��$X)K<b��T�QX4�7��ףV��=~��|��hL>X�FpX?3v'KH'�$�54Xε�;�N^ʿ/hQ�{���I�|�
��?&�� oň�l�Pa�,��la��3(�<AV�� PG:���oz�����H��_�����UFR��l��Y� ���*]�9�Ar~���o3������%w�i�0%�_�(O򬠈��,W��˫F9�4kb��	�nX+�m��LxQ�Dr����3�
�j�G��ǵ�O�2͓��"���r
>>��u��$W;��X6��-{�R��	���H<��@�c5���>�yD�-�sX�1�u�M���j;q2x����C�k�ʥ\!d_ɴ��_�����X���\h��>��[?�/�S����Mp�&��_�)�T���Y�/�*AUt�]��k��S�m�@N��\ܱM<��K�4�&�;f�J/��=e$�C�H���Z>b4Y�0Q��$�h���	e����� m���U^(�)���1U�Fgo�eg�u���"J��e�
�#�ͩ|(�<��dH%{��|nns�}�\6s~�aq��6J�6�[9Am<h�]��)"��}�9Ē�O��:�!���Nk��E6&I(��hF���l*Y�a��,��������9���؝8?���vi,T�pwD~}��H&BO{�19�E�_a�KH�3m(�@R�S��ŁAIb�f�?0�^bx�9��۬钇���LL�(��qJ��ZCG�
*7c�����z����k:r���p�� XfS�~�=X��	)�%��F�t8�ݸjk!��O�|3ۯ��
�#"&$�#�# �{+��(����d�z�{W��$/�Ѿ��T�o��u�D�GӖH��gf��O�m�����V�c�j2#z$���A���~ӽ��
rEpkɻ}�CHiԐC�p�,kd91P��s!h�����>/������\;�z����_�7�z�������q�2o���s�Ē�<g+�6��/��ņ#�c�'��Q�ɟ93T�C�Y`��TTr;���c*9���]���X��i�`G~`�Z����i��!-�Q����lM��Q���x���Ua�'Vd}��Eoy^lK���3�s�k-M�y>�'���c
���;�af�-��a�]<;���Q���DFp3�LdS�_���3�_���BL�^%��ٴ�\�E�n7:W��	CN�^�3�h�"vJ�c�A�����D�4΋�ԍ_8l������8t��@iq
6�yY���M� ��;gx"_gQ�滋=G[_"
�T8 nW]�,OG�(��ᦧ�H$�x~�cek����߮���(�z��l'>T�h�ɲ?,xtrB�op��iY�)�.G�(��܋-v͜,��?�J�{E����5N�]��[�>����3m�s���ON;��V��l����ǿ�G�z�7�������^��!��������N��1q���j�:�jL�����WL�X�E�X�?�� ��O=j��H~@�>ִ���ͅ�ne���2ˎ2dd�NV���$������D�x=P�����A4����t� 2��+��"3�����=�?N�Q3�3�?_�����G!�xz��ߌ��n|N�����{;2���2�)�o!���� ��qr�����	O�g6�>��x7jw�޿N0����ˉy�����۰�������V8�F�̺x�� �>�yn�
Ѡ��y3m�8K{�A9��+f!��0�z����5-�P8R�(�q eo	.����guqGg��QE�j��o\�XG�����e'�&\eV^���m��PJd(_�v����|-��3����y�W���XKE��sb�ɲu"�f(F��Cr����p��E$r���h�v��Or�j5vGj�3�W�DS�?/�Y�;Z��0��h2��W8��?�b���@2�ţ�]c�,j3I����:���(�%Fj��^���C����t�{�9:;����W�P��� ��oU\���,��!�=��aS��P(�j�x]��F��{v��*e�Nu���,*y��cPpw��O��u�;6L�ii�=푷�9���R1V�צ`Oy]
[�xՠ�_� 7�t�+���oea,���%���c;SXio��D>�������{��d'��p�Z>��ޟFb�W�Z�E2�dw�@N�$����m��W�8��3g�`�+?�]<��,���e�7�CD	��)#]1''�2�0,�l{2H���͵�p!O��8z��ʢ�^�s��#�Φaa�	��Hf�����XB��r:@�x�.yS���w�hה9n�Ƚ�٬��V��V`�G���?`(��������rgdZ�ڈMϒU�Y��0e��w1'���B����	*��iU
�'�,e��0���g�-M�O��9�-�3c顃d.�nx�gv�4\"rh����e�ݪ���R2��Vf	;Vs����KJ�#�tD}��uݨݟ���ƶ1ly�^ T0Dڗ����,�蕞���WV�#m�񬂃P��8ת"�	����I R�Ot��-�?��@T�R�6Ww8����\=N�"���jr��kc�R%��|kzc$��^�w�� /���w	���s���	�����ܿ����հ�\�ow0�b����_嵖�B��^}�ٕ�|��-�<r�ͭ�pZ�=��+�]i6j�_�P%�de����8sQ�9����y¿M��M�,�'%�B�3���*)o��I�`������,����L�Xy�^�$�=\R�
�9:�����C���n:6Z-z�)��B����ry6<��"M�]�o�Yħ��T<HQ욖-,߃�����YۈQ�f�Lk�d�h�����s��|�����fE�"�����`�KZ�9��@�b
<�L��&Γ8���9��!���d)Fq8#y� f*�ڮ�.�Wq,�-ύ����wD�t���T9�ɭs۱*C���m1���Yq��o�ۻ�{"=�mV+��'xeO�,w�m/�}�5��|(�/h7�����c~�p��5�(����B�<�a�<���歂���/�h����Nr�N�H �e�g4�E��~�pv��8I��v�Y��S��7�X�X+F���_�*m�
�����/�Ln|/�}�X��J� �愥-R�Bb	V$�����pjB���6�&�Mr�)��.����My�ß�^zݑE�p�;t��;^�85�g#'Q����)�������{�P��%P�����
d�� ��!�d����ym5oq�|��
bID}-n�̀#$�����>>�4�<y&&ͱr�����H2̹A&�k�0{?"����_�jk_�<�l�f�ūtz�P�\W3K��=4�޼�7_+�~�Ld#���xu��-���K�X��h��r6+��q�<�">����:,��}�ढ़W�k*r��|�]1&����4`P��
w�H2�d�X��mm�>��rg�j[�t[��%�?�f��V��>�H-,�:�_�S,Q�.�l�|�4?˕.�E 0v��zD�J߇Wuƿ�vnr��J�DĚ1���ʮ��rgG��afr�����7�ԑ�Bh��2�!���j��Z�j�R�;"������s\��Q��y%��h�*�N蠦sNݛV��1߱n�Х��ȅ��W=ӏA4��[Z�5K�zJ�P���6+p=���?��v����V�L$	�leU-VKφ���~��l2�ׇ�j<�"��5��>����2pXPᅩ��gÁ�)u	g��c&��ۗݍy �`�H�Ļ���U�O4b ��^���f�L�aP��2�Z���6�H,_98�d��1�#.��MfE>SMj��I�#� <�
z�3�DA��}3I�,:Ԕl\e7]��ex�SsM�pq:��݅�6Dg�xV�2ig�L�L�\����8�k�t<X��R�QyN<q΄�h��t�n�.�`A��C+�M:ц���v`���8�����p�2�g��;N�W�9�O���V�pz����ł�Y�h3����5u�f�Hk��/��h��@�R�d���U���ڍ�L��ZbY2� �T)t���(@�J�75��2T�L�]�w"�$M'k��̰9l�GE�����?.�}zN��ݛP�5�/j��\��Ӛ��\�T��G�΋u��&_�#�|�,�٘S�P���"s��G�����@_��4��p�ᰢ^�y�0~�Bu_�Ϳ0M���`y�����<S�k�g�<�lBN��u��^C�F�P ��K��7�dB�\�]�:����ݚ�dX+�m�.�)�'r�U�<�.��<A_�h�]y���\�{�l&��dL��<�̎��=+��ͪHN������7��!�|��&zZ=�f��Ra����$0X�hl�&k�c�g���j�H��\_]���k�%N[cI�o�1A�E���M��L_c�[��v��pI�3"បG�<)��U���6� �%�� oɐe_���/$�
��Vː��DF��w�,=�nJS,2�o>�!K17�5�hb��ߔToX��G2�yEXQW�~q'�#��Փ��̥� "�z����z�1	w��|F�\u� 9��
�.2�I*���۰3d�Dh@�!��.{�iB�	M���Q�/�oc+Ę������mt��^{��8�+*�u�����c@���Nt�l $�%���)#����2�`iT��(���9J|O��R0�K���S�.�m���W�%��zs�����?�ￗ8o���~�FB�@c��r��{$
�P��j<�r�l(�:K+:����U��)�<>eU}������I����x�֔w�8߃�m�I��H���w���m�M����sJQ�;��U�0#���h���@kj�qDB���a�� ,��P;:�m(�Jt,�/����>��v�)K&����,)2e�T��?�P������2��o�<���y��g�D�>�OX��^`*I���S��	'G:����|��I� 
}�'o3�Q����Z��V/�z8�6nm�0��t�n��x%�B��jӡ=ծ`���)��ϲ,�ɶ�t����F��lE��N��t~jö�	�Cq>osK<�҉2��,[��0KJ���Υ|u�Ã��V�-��,~���YQ��U�R���R��$_?����5�����b��"���
ؗ�Z\M�LaB�H�Jݤҕn�����8oy�n8�������E�r7�&*&��lA�<$sd��#�]`*bJ�H�lz�����g�FTn�{���ڴ�*���!��X.����)Ң]J��$|}�JD�:8�lT�3�����|����x�gu�Ù��K�D"�m�2�vK|���ؔ�wxuH/P���sD�SL
'QЯ!���1��4)���˶f>����W��r�;�尿�03�����݉�c�,�k���ze4�6vv�}�C]_QVq�P#�OF�8�T���� �J5�t�3k���ZxP�CC�Ǡ�Qڬ�IV��7�xB*OY�*l�0e����1�D�`��6�������}�э�j�P�����c��,���Bٮש!Y�� )������B���]�K�}���Ix_n�x�������3-E�5L�R�)U�LhI����A1��n�Q��L��_���c��Hjh��
v��x�6ix��GҪC�5�f^Vgw�6�۫T�=�,r�Ӭƻ�S`p���@nS����h`9��������噻�5s�~��\�z���M4S�&��h�I���-4�˕��Kx צѸF��֮��`�v��qDG�(]pR�M�.OѰU\����A�v?}�^���N��v�'�����=� �Qǋ,��gL1����e�
�k ,J3>'Yj�S;�Ow�����7;�5��G1-����,�����WJ�
VK[��s�_It$S��n?d�pT�+���H�l�tc�q��w�݋/�T.Nr.$�`n�'Z�9��̍����]��@`棅�9�Xc��s�.ooA~���@I]��}"+�\N�ڦ�tE����y5�x��Yq}����[r�	�
T��=�Ac���)����Ep0���C�w��Xe��z �p8C�o/�h��ڡtZ�/li`�D3Y�}�e��6c�@�'sJ5��_&N��Ḍ���}���qJ����n���^i'+����b8�O�;��N8Mx�?�{z�ՠk�W0���x���~H�{���%�v6RuYT/DXT���Ձb��,����4L�	�f��n�옣B�'M ��������Q�C�̅�^��u�Vv~|��ɎN^*����(�Ϧ���U,�F[,��~s�V��Q�I�;p�� ��*]L�/�l�!��-�G��ַ�:8R#��w��nZ�j�kT��u�c���)�J�O��יc$*��hiC=�ܤ�
1�RYFS�{��~�+(�GCJ�]GdcU��)�r�$cI��:V�O�r��Sr��W�l�A!b�j��d���1R`�y��7Z��������CPb&ZN���O�}���i�%�=���j�9ф���j�1H�
�U.Ci��F-���_�R�xä����Oj�f�6�m;B�3ӧ$�M��ҳ��i{���'���U*�x��+C3�������^��N��J�Tst2.%�&�A�.��G�@kPI�]�埉������Wy)�|�2�l�x�x(/��&��9�ec^�B9�JX����-h�(��N�z���U��RA �p5�K�{&�i��Kf��[�y(�S̚�X�wSn���Y��,�G-��.��m+��Ё�ð���Pc���b�2x 5>�$���g ��@e$�����������r���Ķ���1AGLDG��4���{�26��K�������*H�n��X|����#�M\�pb<~n7���X�*04g���
����(У5��z2�*��2*q����<Q?�buW-�yi�,����-�LБ�[H������i�����'Ƃe���m�m3#�q�0)|k�o*.i9||?�ȷ(���!��O��!En��T�{�uʨ�b�-���_t {���W����6�̃�
��p��	���"�����1(�楆vܖ�� ��=pM2QW_�"�%�j�%roeV���5M��-�[?���nA��x�;�qL$�7GZ#P�Fd�n�J���8��1�Vȯ��<�ǔʪ�n׽��@�אl����@� r�U�U��)����]�����J�{Y����1;-�FtV���z��~>B19yh/��e������\G:pQ�G"�֊�A��'E\OW�싣�tʨ�i��C��%���g��Xw^$�e�n��(n���5�d��$	�����tD��QEld)r��o 9�GfYx���ُ�;t?FhUc9#w�p �ri��m��G<C�+�l�J/[Ƞ+�/���#�&��z�Z���5Q5��z��3��0W}	���ǿ5��jwgQ3ّN"b5�]��J��J �:�~�"4?)L~��S��M�ڊ."
?�~�NAi��Q��g_a�U_#,!/��r5T��NLծB(�lm�:�[�ں�U�ļj7N�.�����<>GM��ߪ5���f�jT�G���坮bg��ޫ���Y�w��^x������H�� ���1M��Gs�Z��l%�o�'�K�'�[��5�t9�$ӆ��R����c��Ȑ�o��Ȟ�T�k	�`s�����`�����&O�@�����r~b�QG��W�hi�v�6Ea�9���+X�����W +'K��~�^��ݭn��Tm��'+|���V�6��>g�%�\�R��R�sp񇨤� �S\����m?���&�
�'[�:��ڴ����1��C���o�ЎZ+�5[�ئ��M?�L������#K���;�,Ҥv�1 o��q���nvg�bs��ԗG�В��絊� OP�.�P��{��6I|u���a�6�`�a�
��qC$�9p��+k��"@��m�������d�>�����˷�i�&T�
X�h�-9�Ks�8T�kZɃ��j��d@+��|�L!dQN�X���;yC�ϑP�ԑ��i���{�
Zz�g81�&@�@Ý'�(mH�$�"c��
�Hs�����E�TEɫ��k�Tv��^�k����(<�I���3
Φ�e����@e9Z�}ʂ�8L�  Ǻ�#	$�>�Q�#���7xM�{(� rg���J�p�(��J������H�4�kA�lыݝ\�:�⣦]'_Z��,vZ^M7ni��R��^�jPci���
�a]�����g�oA~�b�Wo*��AW���BZ3ΥAb���m!�+DC�H�[n/��dҩ8~L٠m �4ֱ&���>O�]��v�����N�\(��qI\Q1��ɭ�)�!x8� �:��B����Kp	��a���j�\TN��e麁nN+��D���F1Zgw��m��B@И�J��6��N�xn��6�'T�7�/]�Mz��6�e���^Wa�*�2�Q��}Ɗ)�a�.�a�ܠv���#)c��n!ុS3���f/�eS��Q�!Ej}Mp�̛�|�������h�*��JG�䯋\3��6˻GbrD�GP�hЉ�yi�i`p��_�ȁ�ASj���)�co�C�8�|y�kh����*{����̊9Kk���&n*�|��אfF��_M���}e.�0DԪѫ��o�D ��>5��Ȓ���sɒF�&R>��e�����pѭ��v�0�:�����:�����m2������( �(�j*�yn����~�j~b��ʈ��zǹ�plb;:��?yg�	��ζ���u����|"?�!X{h|D|*���K�Al�1��WE_���*t�����{�B�8��^��
F��'W�ё��q�q��+ƍCQ�}��iL.�*,ǻ��S����gϫE�.3"<���]��5j\n�]r��c7��V��m|pd��H��3gF]$֊C<<q�
:⌞ҋ��^QX�c����#U�x������bf /�҆{�/��Q-}nL�Ok5[S	g4�]��`��PQqr{�fO�J�Ll�j��K��kuJMy_���Ajj����&�~��c6e��QK�hť�*\^$���(�]��������e�%�W����f���(�'��Η�R�z�~q��¨�F���o���}��٫���}�|IV����MQ9��T/�B/5�jk@O9 W�TD;�e��y�=��Gh��޳�5b̉���9�t`<7��&�/���N�@�M��0��<�Jl=`�ކ��C���3���K.[d&)�9��nwJ[З*�OǸn���D\̗��ͥ�\tP�h�vuU_F@z^�����������P9��Q՘1;JQ�tN��9z�U�@��w���3���2a����)�>�3���{����ih]���}IYM�Z���B3Y�Ӡ�λ4 �x,8�&f�-�+%xV�.R٘�1�n��t�g���
 2�Mx�G�ɫ�T%.A9&����V;��vO�/�pU�Ε01���I�E��Z�ţd=<���!���� �¡U�x�g�d�y^���(rXj26� BW���)�����Mn2�h���XV�o��X����>�V�)�,W��8*#��T���z赈�}���6Z�iiU�U��i.Y?g���LZ,=1^����x�)Io<�]���V�O2z�1:U�V-��8;[{Hջk:[I}�&���2��7lc�]���D�����j���Eӹȩ"+e|aLo<t���yz���l�Ͷ~0S�!��%"w����-/�RL$2,�]�{ӟ�v���!��j�A/���>�X�����r��߅b���;!aש�J�/�n�<^Z%T\�����ǀVtΈ���ܳ�&&������s*���&�s^P�1i/0�=;���n�Z4�h��`t~3��';Ⱥ���L0d�6��U��b��>�W�a�����w'�l�=��#:BP߿���X>��XS���4�s��M��U4�� �ɋ�:�����ԡз��3_��sb=X����K�j?�ϩ�g�:��%fR�* kIw�x�y7��B<�G��ʀ�kj�Z	�q�ֽN��'ya�퍻�Um���ә���o��ra�|�(�q�(�b.>�IIb�eɇP�]}����{�� B��O�38À;}W
��� 	Sg]Dd�[��]���fSʎ�=��Ԫ�:G�j8��C��)H�������4Pdza)`K/E�!�u�z�5?K�~j��(Y��+��R��� ��IQ�,��n#��r"��JXm�H���Q�������$�%�����:%pTKAG�����	ek��B��:���M	el3�����؛?�:d�Ɗ�L'W!�C]����q)��{iuQ���4�wLQ��2�mT�	�c�0k'��on�<e��-��=��@�q�F�})���f���Z�`���}?������@㽶]�e4�-{�,5lb�jU��D� LrJ�ּEs�8�wBo݊��tW�Wwl����P��r����p/�F��O���\x���6Mbwl�.D4�z��>�\�Z�Q>{��.��9NQ2-�4Q��ZA��ƈ��b
���b/
W�\�0X~�5���!m���Ļ�\���|�=ՙ��n�
�x�gaVm�~��������-�]�w�x
�s�z1��;�5t%�V�0�ۗ��W۔i*琬�f�6=O��>�^��[������B6�& �`���#�={��_[(�vJ� �py���� 6����e��A��~�P�7Y	���G�("�i�d1�	R}0���9O��{,�׋����]�+-�])�=U���5�Zf�������K���3�7R�,�N��|� .z�1������	������{���^��tH�9���D|2��gf7�݆ʯ@� G߲(��Jy&�a$4�L<��Xk�v��C��R�C���7���,�t>��̭���jQjYMda&��yt�����Sl<��2KF��͚���Ňd�nү�o${T����n�o�=SC��r�5v�h��1�`M/ip�g@Uɠ��UK����X��ӿ*��\JR������c@_3K���u�ɏ�n,�e 1���?�$@�ڂ�TtWX��)
�o��h��Y��p��b�����E8�蚼��W��N�iC؛p�*���tUteKϼ�*���*Ұ&<vɴ<��a/���M���̬=�|-�!ՏC)WD���!���uQ]��7��E�XЇ��l���T��j�(�,|�8�Va����o��O���^(�@���W�q�O��*]
�ͯ�O��@o�
emk��k�j͂�DI
rs�r�T�����4��^]�r#��.��wz�뚧3�zSJ�������`!�c���b)q����F�)v)-�½a���ޏ7S
��'��H��V0G�3g��]7����������V��\Lb��5f��(@�
�%�fG�������4p�!��1�Q��ܕ[�7�x;{�Ӛ ��0A+����$VO� ,�x��́���uQ#@����ᘹ�3�_�gc��'"��+�����}��C�dRE��Ϸ��צ�FR���j7����Qa��^꧐�Q��,�B��FÁKb�xR�/<~�5��]ƭ�p�9e�M��2�\:�o�c�z����ȅ[Buq��.V�h�bF�R��Q�l��;;>����V������d�����c��G���xpMipY�DH���ޡ�OI����_�F|�ni:04E��T",���A�T��V�&0s� �m����c��8���{�,�h`���|��px�m ��/d!s$�ϑ�˛�xV8-J��V��S5����VW �ݻn�U��q�N��?��<X�d謏�"1$�%YA0p���d>קAlޓuz�d��ڬP(rdf���-��Yʃ�Y{=�*H�YD�AL�z��=�LPE��M�%~z]Z���#��,(��"��q�Q����A���\���cߜ܁�A(;u��Ü��w�_kLܠ��S�=�뷖L�ذ�췠���a_�̏;YK�Q�Z���~q��w���*�h�
�%���u��*.w�sp�+�#����2�V���1-2�ɯV�Z^q>qO�щ�CUA��!�}�S���Rr
/�2�t'�����{N�,K�pj��tt��2�������=�t��)��1�h{�y<S/�&���|��()Y3�V_7lUh���Tŉ�8����;��A�V"
�z�ˤf����N<إC`tF襺�ӛ��k���
�*����\�Ub��	���)��5����C\��,#�]O[��71c����F����B���é
�Fr ��N����Zh~�;t\�{b��� �H�3�Xn��J��'���~Z>�OJ""��ȊF�U"�D{�0�*_�mL�y�,�-w�Gzg�r��=S��[bTM�>&�/f���@���	0ILkn��VR?�-�iJ(��˼�$��Z�̽STh!�ǥF�=�A*Vl^l.��m��u����Q�Y?
�Bi
�e�?���fh��|��uD���աZ��R9�k��-���v���4@���{8�I
�F^��x-�%+����8 \!jSH��A3��,�XorV޻��:����x�g>*fd��<铛�D�47�:�oS׷�"K~���q]좸�g��^�g�Ԗ�A"��ZH�t�|����z�,z�a�s��в���ʇ숝E��^�a'����J:�VI��q�#�]#b'��8Yf��rr<84Z�B����q���f�:`7$xIeο��d������XY�ƂZc�Z���-3���jV����/�`�$����t݀�6�cքP�?��U(��May흎~	{J��]~)�(�%&��Iz<��o�m�y��klY�qYR��y����A
��'�gN(������)a����CǇ]/Za>�e��a>�!��@3�qs"}����<�`�:ռS��W���Z|�ʧ���)�|�t�M��������[@�IO�emue�Rw�)�$|z�DSR�â45���pxv-�er҃RIb�} �:� �*�+(Bg�L�����$i�B�MA�@����k���/���s'&�o�����Ժ�4��r<D��9��j錖(u�=�	��
�2�ԒGhTs�JVTe�w�Va��:�0����cɲ|��	�r�����Ȏ��l��:	\m	؜�g��x7�%�f(�`�����47r�@���I
7!�1��� ��3p����<�%n~��I�J����=�� �@`.P�R�2q���"�{G	+�u&�xSxm;�S<�Vߌp�l"PR���1u������g�7+��.ck%����J���S��F����UEh����a�Om;�N��s~����W�7�R��K0�lAx,~n����t��=���Ƀj����V�:�$�j�uk��'���a�q̮R�� X� �2���! W��K3�Lf��@�Q��mC����6�p�Ң�?;VK�"�V*�`;�,$s"�U)�#Q�Q@��q���34�P=��K�q�S8I0�0?dN�Z	��EV��I�!�i����{�5]��倝��b�?��Pٚ	_�V����j�K�O6�3�w��p��{NY'�=�J� g�+��z}&&{�����jTm��&H�+��U�;%6y.�zX�V�F#�O�5�1$ŷ'<lbk*�@z�J������D�|:WeVj83�n����"��'f�Mr 7�1c,�d�� ������0G������v�+rd���S�U��U`$kV��J"<t�h}�����/3cR�p8�uUx��Ȯ2�/�n�X�K�B7����Ȑ�X�{E�Υ�����|��Q��b�V��к;�������
,"�Ƌ�s������鑣��̪m��E�Hв6ؚ��\{�MHժB����P�=_��+f|ӹ,�Bm���Fm���9�
e�K!��{c(�(�h\7R���������wꍒ(_v��	�yGɁ�cR,c�"��)vK��m�8�۾�^�����w=դ�A��90���a_���`c�U�mqz���������������?l�{z�U?�'��pX� ��O��>\�J���~p;V��N��(��t"�\��W�s<��4��	㕦����
{�WO3w�s�ea�8�Ѿ��G���8q�l�#�7�����c�	[�$\7�T��1�$ݥi��(\H�%p��	��Gk��<yq
��A	5����d�w��ŅM��Z���Hٽ@�Zq���K�F�.��`��qu����:�˧�z���ehN%�L�ia���e�OaP{"p�'���V���v3̶�mx`�L��k`�βkn-��S�J�@��k��[ֽ��UL'�����z��m
[�w�i{��-���WoCH'��Y��H��c���Ar�f���о��Ab�L$�F=�5
��@��S<����6�%��$��o�,�R�N�N�
�,|��{���4u�J}�}�11������}���