��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$��7�4��L+Q���+2�"H�������v�ao4��	�u��=��d=�>�iV�f��l0�Zs��7���~rM��U�`���e����K%�u��ݒ-� rā�SZ )����C.��&0C]�-��[�3�-���+��պݣ�k�J�vo`�A�����f����u�X���v�=�а���]Q�Wۿ�߸�=_Q�X����j>��Zw�K��SvX��ƥ.���#�����Z�0���#7{��\S$��@1I�QX~TQ�E��db����۰� ���>0�%�9�j汈��}��1� ��2���h�G��SeY�a���	'<x�p��k�H`�H�j^y�0�s�78+���ֳ�`�R3dW��_��{p[�?$�s0��#�zS�_��bH
�c�p�IL7]� |����Q�� ��Rr���=��E즕2%�����`�^��l�q-�]�p��jf��Ӽ-f%H���ȳ�>��+���M�71��4_�) 3�46h�rb�J�W� k�h~K0�>P$�_n)���5�r�j��W�J&޴o��$>��6��ŀ�;A~<6P��K�~��f��*I
�Z��}`q���ApC��n���g���3��-�іrO�mF���,�$��@�BI�q�}��Ȥ֐����î�䂧��@������U���vU������ �T#K@f�㯁����|95<@���+�-�)�����K���FI�k���*@�m&���
���ma1[�2�u�I�\�U�yu���o�|��2����;�W�W�}P�K>%5�'�8���׫=����k��,�t�M�0�8]q3���N���GvZ�i�+ C�e
��Ќ�S�v<%���q��e_��
�k�夞��>ZO7E~��5k�TW Aod��eE���G���ɑ-'���?�G$����ќ����8ɸ+ 5ʗ���l�d��,�J�
�^�3b,�����J����#n�zK����z�&��;|�\�^���'e�W�����">�w*<���=�O�V������0g�R��6�a���=y`(�$g�?���x��L��䧨ʴ��<�6�}���0�&�IX�b����#����g�ƭ��wކ�C�n�n2�1�N��0�Ã�ă|Z�k;�&�f�(6�7���3�u�����P��3��	�ǝ(��p��)���Sf��l�(��CIn*EJHe�
�*רT`�a�T����|�U�����r�����P���\o���G�j|x\����<0?OȾv���'�?h�>��n1��Im7�<�Y�vΔf�U�1��q�֢�,d��G���X�^����8|HpL��T��'�$6*��q����
G�G�X<�@7��]'�̍�G�^`,4��In���4azl���<�z�D� ��{,�A_�ّ���|3:p���wa�C�=wd��74thi0�T{���>Q9�JMG6�Y�/7����@����i����ݚ���v�Pű�R���nY�ī`u�x-��
�+�U�0���s&�Z�W"�xf�T�^b��n����?\a�y\�=�V�3`% ���رfh�F��rF@^o*�@��M�ж&��%��-������w��2y�C Y�ȶ����~W���}GmW�����ŉ�ϣ(�PKz�8�v�Y(j���(��t6 ���\R�n�"�,�u�@�[ڀx㼾4cH3��&9��
�[�]��������cphY�����b��=�ch$���;c����|�6�O=������x�!���
?~��7\Ԗfi�(�gZ���4��u^�w��<a��'��Mzh��ַ�JW���QY�gce2�#v<�{*��tNo	8�T�����O��n-�c����'GYf_VK7Ǌr�@?�`	_!���EW����Z߻)	3k�,d���|��/�\83!�!uY���ڿ�:B����#->��7�m-�sBן�e��N�]S����ɏu�e��wL�'[��EZ�ܻ�E`'�0�_�,-����tx�[2p7�\"2�	g����Bg�v;Rg�Oܔ�IJPW \j��ѷf+:Q�w*�4/��ە7���K�]V�O0\�� P��肵�B@u:�^h�`�w4�⺠Y�p���a�F��14�(�7�T3]ԖeId�%{b�u�4��*[|�Ȍ㌡��GF�a`,��Vu&2�l:#�a��B���Ǵ��G��?��Uh�R���I��7�uS s�rQ�2#�n9ގ�0&�э�)�Ul}j��{U���N'�[�b��#ݐUoV&g�3W`ނkK��>���� ��L���q�ָ�$��Ų���|�-\C�?�S���ߥ��e��#.7ϛ~n��~P���%��W�It ��6�u�14���%�16���6���\�3�"L���76�����\��Ɛ��R`TvP��\�>٘�4d4$�&-��V��%왰�9�g �k�#7>� �\`	z!r;�vL�n�h˖�����Qٺ���ۑ���ݿ��o�9½�v`P�H�al>���9��d�������|If�)2��Ml�y�qg��z�j�p����c���X�;X�DM|�&������~��D�7��WHV�.�h�I;V�T��L�&����c�2�%��&:'��yw͸�z�5��Bvӯ��qvL �(��a��_ZIۛ�e�,�{}�!�e�6PZw��+��)���_�a-c��ܡrV^Ubd�)��@~�]����XJk��>���*�r\��DV���\��*
FbZi}Z���\�"�[9�(5�J��5|��VA������<6�\v��I�̟����A�!���!핀�i�E|Π�� ��β%eF\_,˿СG~PST�D@�.p��Or������P!�z��_i����)n; �c��o���kZ�M\��>�3�{�g9��A��oV<C��{�P{����������&T�����V=&Q0W�=�1z?~l��5$,�}�P(y��a���d[��ŷ��}�H"���L��&1h@A�'��
�!��}A!�*�Fe���\�_T�37�2�9�s��$�6�&��(_�-�jYmG��D��K=n�x�$�p�po��j݆���@b��݊��L�ƭ�*GZ~w���wbe	0e��Q� ����5����Gܞ{?L^ � 8�rx*bN�V�ia�>Z�O�찗��t���E^]g�,�1y�Í������U[P�"v�r�q{�� s��B@���PN)�Rˑ!|�`#H��xN��t"q�Ӹ����]b��7`�ћp��7����o���w�?��GOߴ̥�