��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� rā�SZ )����C.��&0C]�-��[�3�-���+��պݣ�k�J�vo`�A�����f����u�X���v�=�а���]Q�Wۿ�߸�=_Q�X����j>��Zw�K��SvX��ƥ.���#�����Z�0���#7{��\S$��@1I�QX~TQ�E��db����۰� ���>0�%�9�j汈��}��1� ��2���h�G��SeY�a���	'<x�p��k�H`�H�j^y�0�s�78+���ֳ�`�R3dW��_��{p[�?$�s0��#�zS�_��bH
�c�p�IL7]� |����Q�� ��Rr���=��E즕2%�����`�^��l�q-�]�p��jf��Ӽ-f%H���ȳ�>��+���M�71��4_�) 3�46h�rb�J�W� k�h~K0�>P$�_n)���5�r�j��W�J&޴o��$>��6��ŀ�;A~<6P��K�~��f��*I
�Z��}`q���ApC��n���g���3��-�іrO�mF���,�$��@�BI�q�}��Ȥ֐����î�䂧��@������U���vU������ �T#K@f�㯁����|95<@���+�-�)�����K���FI�k���*@�m&���
���ma1[�2�u�I�\�U�yu���o�|��2����;�W�W�}P�K>%5�'�8���׫=����k��,�t�M�0�8]q3���N�u��j�������ZJy�H�[`���W��b���-qJ��E����5q\bx�w>Ʀ��Ò���r�܂��%,��HഈdV�A^��k���ɖz�@�����K9w�5�i~���^��V���.���v핣����KXb��gt �K�1�<G��R�2�Yj�܃�)��T8յ�}𨁥�²� �r&�S��0O���d�kW��;gJ�7���� P4�ꌄ�F��0^��@�ҡa3y����KVS�E/Mֹ �.g�Y�;O5|B���9��d����av�VkG���<��-�KȱFG(�=NI��N����Ka��"h�)^�e�6)H-�{4�e{=p�@�[q�S��p�Jc�������N�o����"k�!�J�W����:he�
Z�k��6�>U0L�DǏwQdk�Pv7��N�\�1�Xh�	C��X#����S}�K��{P	�w�d���[�8ǎ�圊ԓ�R��sX=��-�^��@O꓿�fhC��o��䄳��4:���q�
U]�kB�̺���	Э���=�ŷl�X� ��t/��?~�&��[-_-�n>I!H����꿟����Q_�'�ܥHN�C|�o`�#7��m�.D�r��)����y;��Eh�>3���~N�X���8�h�>-���j����~,��sx�Hb�rdQ-A���o>[v�8��KF�B�]KB�!
'a)D�G'1=�	 u�`����Q8}�����y���N�Y�C�{�w ^M�c��V�����r2ױ���iEI�m �9�	�����pN38z��� j_r7푎�{�R�W�^ ��;���ky���_T��x�r�����,�
���圁��qoM��s�Q-���M�Jo|�q��!���,���[�d}c�u���u�O):`s�:9�����'���m(�P���įQ�fUB��ʊ�U�Ö=�����5Ӂޏ�� eO\šR	��+|Rn��B����B8�}D��M�J8�I�#�/�X�� @�����od�������Ag����ȅK@8T�v��t&vtr��z���?wd���wF��B�yv�l> �h�Щ
9��Y�x���\SD@,�R{�3��:
���\�K��'����:�V8��.��|{Q~/�e_I#r�.�C��	m̦KV����3\�1yZ5Q�=s)/|�����P��Z|E:g�q���0y�J��� �΍	m�If�k�0� �x�^T��K��Y J��aS�T�����І�V��u��ߛvnM��j�x�!d�$K�jT}������d����Oc����3�>%��6X`z�]$F��*(��9��J-�^�����(�����69��"2 ��6���P� ����=�gmy@]�oW�f�ⵦX?�������0:Ә���҃'I��������{���Jm�b �@�oe��etw��1�!�	��/A�=���.'ma<�+�.�a��[�2��_���!��m�A��0M	=%aA��t.�eWd��� ů�w8�bk2�rV��9�}�Y��L	[�9L��"�˨���8���v���7z��j�a�SI�n�6ȍh�P�G��*�5]�b���Y>�r�K��[غ7l0D�՜�J#i��Kˉ�mqB�N�}oU�-5�h�1�R�9/-��ws^��\�Eg�,��j��������Oy�)���v�W4��'a#\ֵr�z��
���;g5�ɯ(ATߚ#ffGVB�Y8��!j�����LP�sq�y[0��>�>���Ϻ�*ү����9g�|��D�m��K��b�e�ԯ�1H��P��␱�fgȦX[��/f�
�գ�/�Kj^YH���f9ʣ.��0T�q�gK�DOS��So7��o�"8�i���K�P=���"Qkr۹�'g��1�d��&6`�|Ȫ<\�TX����.z�_#���"�����a���o���x�XUXk���t��"Р��Zȼ�Ζ���J���X?��y���^����7��g��E8۰�*�"8 �]&���
�l�v�g ����
�g�;�PgHM�$](/�������w}?:��F"��ս<��qQ�k?-ߣm~Z��j@I�zc�%�$�4�Pmz	�W�������l�>�կ��:� gFO-��'�0U�H,<��$����ܺ��N�+��,���'�|�������C���/��7\�BZ��A�|���-���ޫ�Ĝ���ԃ�N��"��'� ��-�2p�)0~��������*��	?&I�	n�+c�a��(��V�-q�Ғs@le5��hgk_�N���L׮=�z3�w�]
 �Mo���ߓ�e-��gS��=�36��e����R�x�ʟ��z\��M�rfiN�~7v�XlL����QoJ�P2��C�v�xN�:=o~�:=Rmt]���c��5�~��oa�r�l��2f��V����Q���RJ�c4��׆	��E�[ۥ��.�s��VO�.Ҝ!̐G's�I�͊;���B������QEd�.���(���F�Z�ź1��o��Y``y�
eB�JH$oڈH�W_���߬w廒�2l5E�eLo]Q��W2:�*���R��9��
�^N����F�f�4�9��sȐrwa�pr�A��J��@�;�����4�4x��ρ0����� 7���4��!��=�31�JZi�[��p��2��i�o��
�t�B̮zb�PL��jð�ـ��mtr�g7�ֺ����^dm�����\%���1�=v��mqdT���g�Y�
A��Z\[ć0 
�������U]�~$@R�U#�A�)��X��9�Z���1�����8=�-��U���[*�����ܵ�2Toݦ�6����_���"�3����>��<�u8�l�Y���%�</3)C,��!�9�7�|  �_��n̚�,H�A}o�V�G���.Um���o�<��7�՝ܴc����ON,J`�Vf���C $F�_F�#�*D�Ԛ��E�j�˾"@3O�u�0Z���;�{y�
"^d�o���{�F!���Ҙ�=���6�SP�<�
�q��/Q�"�o$�$_059�����^Vi��B��	F�Ik��������wFqV�F�Map�А���4P��"���)G�zv�0[��8Bt0�R��JNXStR�@_��\�S���I�)�۔f$��������н�l!���S\(����G�m8���Mys�'@t2�6�;��cH"����BuN�5�$N�3�^G��B���0��r�x�����/,�l^����+��24f
)�#�:�,^_�yR�^�_iz���N������Q�:*��"�	��_馍N��<'�أ�䒰��J56��²<����%�����d�zV�hg�K�#�6��`��XQ��������C6�ؖNm��y
�	!�'�6V�"d��� by(�7�ɐg�42�Ⱥ|&��;�H �f��m����D�|@��skԏ�7��E���$������%����yJ���[Q-���wfs�	�]5�bzLV��*�7l�[,X�ܑQ�]~5y,B�V��z��.UDZ4��D��=$���nK0��E?���0]TV�`|��h��;%CY��Щ�_?P �Q/b͔a��� $A+2�u�+�/�:lڈ�Ѿb�0�����Ç�`
:ξ�7
�J�˽M�Z�ΞX
�9�D�}�V�5�Sv"�B`�M̙�Q,Zu���߃���i=�zXARw��$�N�r ����?�ח�c��q�F��b.�Rn>m)�[�E_��ev%�ò�Oѳ�r��Z�7�Ҡ���S��i+nrYN�3�hN�"���ua��v�\ݺA>��l���4����r�?�P<�wnh9pΌ]���F�1�6J¡;:� �ұ�/~)��5�D�W���u�r�Htt_^?�Yy	��G$��̊�~�Bk��J2I�Y�0���.�ܮ���)t��U�4�Q�W�	ô�+裼)g>u�Hvj���3��铡�������{fu�� 
���H�K����g����p�����L��]J�����u�-�xC�b���nȖ�eS�1V�96��y���)K�;�YI&.5(c l,�o��Fyd���_,�?p]�<��)g����l�?�w�67����	�F��� mL~��3V���8����?k<��:�(5��O'\���^w��"J�O�%MyEu�I8k��n�~�l�!�(�\~�9/QI��y�9 |���]8с��+�ɠȁ.D���t߼~�T��D�SyI��N��Jm�)߳J3�F��EƐ���xO��F\d4�*uV`4_�z9��A��bZ~ �d��s��h�;�]9�o�(��,����$��E��A9d���_��F�����MB�Ƒqp��
h��x�Ykʃ�(�O�'/�[�x�Pc�bU��>G$b�Z�D�C�AⳋB
LG�c�JIW����+��"�Y��Dd�!�cMd�Q����5�J�}�5��F�Y�6]χӲx���\`Dc�{f|Ɲyf�~)U��X\$�s�����zM���4���Vb�ha��o��8���(��2�+�Ė@�f�%�М���ܖ��&5��e���C�k[�|�
���̛��H#I���Q䰊P#SEs��_�'2�){x2
S��<=2�N���ҏ�!��w��#ܱl��N��p6!3����] Nϐnvb�H�8�Mu�i���&���~
�|fJ1�%"����4�x,�o��o���n��/��F�F�oEJ�A�$�*�
K�b��zՌ�ǖ�4g��8C�3Dry���f���N��4�B��}��T�,��w��DL�x�q�`o��Ǫ�7��#f�J1����aW
3���Ö�;<+�^����RT�e@����x����Qx ��z4F^ָO窾݃���/-"Aq�h���Wo�B��������I�0JԷJOPL���6���)�g��"�«u��Qvu��x�Ӑ.t�^�=6���k�$�僋a)��V��'�� ���.��zQ��<g��r��d�+l{�t�S� *�0o��P�E�ǵv:�F���"��N�7�l"��܄��y�!�;�'�rI-Mm_�E�ªJP���YE7c����cV˳/3_�B`?�G�q_q`akw=�7�/+| 0T�f겆���pA�R&�&�^�m�
���