��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� rā�SZ )����C.��&0C]�-��[�3�-���+��պݣ�k�J�vo`�A�����f����u�X���v�=�а���]Q�Wۿ�߸�=_Q�X����j>��Zw�K��SvX��ƥ.���#�����Z�0���#7{��\S$��@1I�QX~TQ�E��db����۰� ���>0�%�9�j汈��}��1� ��2���h�G��SeY�a���	'<x�p��k�H`�H�j^y�0�s�78+���ֳ�`�R3dW��_��{p[�?$�s0��#�zS�_��bH
�c�p�IL7]� |����Q�� ��Rr���=��E즕2%�����`�^��l�q-�]�p��jf��Ӽ-f%H���ȳ�>��+���M�71��4_�) 3�46h�rb�J�W� k�h~K0�>P$�_n)���5�r�j��W�J&޴o��$>��6��ŀ�;A~<6P��K�~��f��*I
�Z��}`q���ApC��n���g���3��-�іrO�mF���,�$��@�BI�q�}��Ȥ֐����î�䂧��@������U���vU������ �T#K@f�㯁����|95<@���+�-�)�����K���FI�k���*@�m&���
���ma1[�2�u�I�\�U�yu���o�|��2����;�W�W�}P�K>%5�'�8���׫=����k��,�t�M�0�8]q3���N��2�P��@ۻT)��8A�G�Wc��'�-�B��雎��C<K���"�c
�@�J/74�?K �l�q��;˝(+�����.l�2��ֹ)�wC�8o4&��3�C�5���-Am~����u�bX��V��$'��5Ze�ǌxz��B��M�-������d޼=�{�4d)���T���Z.: 4
%k|w�0<

�ƛ��+eWd��#M�Н��M;�/�����<�yt������e��&���mP{���v�Y�;p����'*��gNG��|uǗ	�^��\>�gUJ�Sfo�� -G��fI���99<��i�s�P��ӎ	�4�J}�L�L���%�2>W-.E�b�̫�7����?�H�0��#�ut_��l�~���v��/�R���������-q�S��T��(8��
���7�0>G���| ��/��*@y�����'��$Qn(�t!�44�MA��|�=�.m��g<�l&�`����W�G�f��T������ё%��ż��n�G2�t��`�}y�9��	�c8�-%����Uĭ���]��`TO�ME����?�֋��|�`�3�D��H�l�]���[�/�E�~vLF6xq}�a.7M,p�����V�^��_�l���׌Di��j�+�fg1�tTr�c��^��e3J�Y�m��c�d�ُ��p�Q��Σ�2c�	muQ�B�҃�N���5ܽuJ8��n�&!�L�*]Q�e����ʇ� ��)�޶x)A�\������V�l��v?�j&�3W���8�VP0 o�j�O4��w�*T	��X���h	�AVeFI%?���M�-����$