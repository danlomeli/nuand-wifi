��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� rā�SZ )����C.��&0C]�-��[�3�-���+��պݣ�k�J�vo`�A�����f����u�X���v�=�а���]Q�Wۿ�߸�=_Q�X����j>��Zw�K��SvX��ƥ.���#�����Z�0���#7{��\S$��@1I�QX~TQ�E��db����۰� ���>0�%�9�j汈��}��1� ��2���h�G��SeY�a���	'<x�p��k�H`�H�j^y�0�s�78+���ֳ�`�R3dW��_��{p[�?$�s0��#�zS�_��bH
�c�p�IL7]� |����Q�� ��Rr���=��E즕2%�����`�^��l�q-�]�p��jf��Ӽ-f%H���ȳ�>��+���M�71��4_�) 3�46h�rb�J�W� k�h~K0�>P$�_n)���5�r�j��W�J&޴o��$>��6��ŀ�;A~<6P��K�~��f��*I
�Z��}`q���ApC��n���g���3��-�іrO�mF���,�$��@�BI�q�}��Ȥ֐����î�䂧��@������U���vU������ �T#K@f�㯁����|95<@���+�-�)�����K���FI�k���*@�m&���
���ma1[�2�u�I�\�U�yu���o�|��2����;�W�W�}P�K>%5�'�8���׫=����k��,�t�M�0�8]q3���N���GvZ�i�+ C�e
��Ќ�S�v<%���q��e_��
�k�夞��>ZO7E~��5k�TW Aod��eE���G���ɑ-'���?�G$����ќ����8ɸ+ 5ʗ���l�d��,�J�
�^�3b,�����J����#n�zK����z�&��;|�\�^���'e�W�����">�w*	FO�Δ��v���I�h���/�*n
� �,�/�����3��� �bт�%��r@�;����s��n�
e�%!
P�'�,k��
j��l�o�[5�+�g�B��cI���Y�m��dU3��&���Y��3.1h�������t���^�'����O�D�F��B��~'DT��[(��Nˁ��>$�Vv9c`T��;[����d�$j�a����{�׫��A�vX��G��\��ܛ��Cƪ JLNb��&�L:42.�S����ݽ��7�3	&V�A�XIJ�o흕�p����t߷���]�����ڑ8���lq�m�Y�p�?�O������p;�	�a��*G�z������p��b�4#�%\@�˖dK��`��3֧䑛n�TR
��d
7��G�w�՘
ګ�1��1����b�7�y<IZ.� g��"�g�7=>���!�rx����;�����,��G�ˏ�K�9�J$	�e&h��j��cţ�w����QN[�R(k�6Ӛڏ*���DZ��K �<H��3��V�j/ֻ�ظ1���-wy��[�f��3g�� 
�3�E���ذ�A�s� �x������m�$r�e�O���N\��d���SE{A\�B��j��+H@�E_s�(��M��x�ǫ�����-v����y��篼K�-:��C?���wi��Ժÿ�S��]70����7�.�E��9�������&�֖1�b�Y�N�4TS5
Uؗ�m��r�%��������$(ov�3{_F-O�u�X�.�� �˃��y�V�/k��J�P$ef�S����*K���;�<T��lO�)&��G���s(�eB�S[�m�x���Sf@��L����`��-A��"'�H_��5�� j#
���n�q�E��l����Zi�d57�}�J�R���	�ɾRr�D3����
�������TݻY�j;*��L�e�S��C8P�AC��f���Q7�	i�;	�u4{]��2�*��g���_=$=�� �u����ۏ|�$�3������(˘<U<_���/	�n�p�<p��%G�)~������m�4K�(�$�TNGV�o�,��\��8� ��������i��ZV�`s�t�ȩ�I���j3��q���?���q8^^R}z�X�i�/�͍�G�qʟ�-��(fh�!��Ʌ g�gA&7Ip�L��U��<�`<!�M��L�>�h�<tT�e�Ӗȕr�_S�����d��r�F������X�H�k<�Cݒ����s�C%=sP<^����&5h�RB��gڸg� �29Xq�K�	8^�R�{B���gw_����,.AW#�^����SR��^V�`W��Y% }#��݋L(�m?pݑQ)�)�E\dsI
=.?q������8��ٷ 0�{��a|�뼆#���o�h(�MU�6r#���e���/?Ӭv�����2e$�u�Þ���B��'Qt���JN��.蛖Z��8�C����	w�0��-�b�ԋ}|x�y��0J"P�'��2*:����?~�ck�T�Y���L��#��	ld�4��YY/yu�$��ɖKF�w�񵕨lrV�x[t�a�f����&b�C ���c����|P��C��?+\�����:�>�ҪK4��Z�п��AD^�w3�;9۞�EwJ��F��Y@��ϊ�×��4#ײov������F��ؾ�e�v��,���r�v�Fg�OkXޓ�'�)4����8��	�ѕu�29���O݄�g�>݅�a)ʕ��dHn+��ױqq���~7��9I��)�SꛢW����sy+�d�63��:b��[�9����bn;slzԵ�6��ʩ�-���C��IT�Ʋ���j1��h��]����t�w�QC�-|���h.��p](~��
��̓ʐ��'?��P[y��M�/̤�ă)Nt�	���~?"��wp�s���?>��>T��~������#�Fx8��#�?�R�V5���^.�|�a������`2ƌ�� ��1���/�x�J��M`����:��~_Ћ-W��O�3g�+����lwCn������Օx�hv���l�VK0����+3Qt=c���Bt��tZ�@D��i��$+��F�0�3�^�M6:�۲B�K����F�ԕ�|Z�L�N,�x�#@Ƌ����ˎ��/H�>.f�{�Y��*gX��cR���/l����S�� �|�h�P|r(:���+ōw�d)���iW?�@�8��JLc��O7��H9��0Rz� ?A��sh@aM�Gպ�ُʲ
�v��m��]F�Ʈ Vc��.���/h��US��\n�Y��WG,��SB��	gdy�:zq%�eO�c�NM)p�����>8I �UQ�W����6��L~�<~"Ĝ*����`��2��(��_S|�ED�JmZ�	�<�D�y'�#��Tw��:Ϸt���^O3&�m:3ȟQ��m�����9�KqG^�cJ����a���g��V�2ܴG[����_8�� �B�߁=/�����X^큩���Ǔ��*ȝ3)�m��t�u��k�qJ�6�~��3(�"�m�K��E j�Ľ!6�7r�SG`Npz�����tj�L�X�NI�L���n��0s�}�� c��(��u� �<D��8��u���BՒ��l�[Wi)n��H.�8�ֱ6�?���n���=Kڗ佷Lf�dӿ���DJ�7QlתYC^��Ru^��H+4Y�X�/g�.�F)�$g|*� �H)�t'��R6����fi�խ�U(�+��0�2V\ɺ�h�\n[�H�.i5��T9��"��d��Y��P��#N���o����V�����������y��Bݟ��X��A��U�qN�)��7F�����!�w�ܗv'���M8׆��x�&9���r����;=A�Ǹmq��f�Lќ:��o��m��x�.5���ns�2��D������;�;͚@i��[y^�B����Ǹ �8�����8�z��l�$/+�hu����U�	ù��6 5��R4G녁*<�N0䣳8������$�z}TM��-Q�2c�����M}�\�׉� ����=k|r5X�*�%���[f��U{s;�
	���ne#	$���%��7}L&�6S KjK^�z��<0���p�ّO��ŞT����^�M�f��'l���̮yI�?��P��Ah�����N�l)��.$�:�Z�nE6aJ�2�o-���:;��1v�-A� �'2� '�����0f"��/�q}k�9�<���ߴZ.Hj[+X~C�3�p�7m�ja%�xe�M'ψB�^�w�ʵܠ
��%@>Q�f]	J��JD���Vj�GNz0:*x-�bf�:hMm��ix�R�Q(�>*7�t!.�.��~n�bg�b�T���A��/�*��7`A��.�T�,���s����������c��0 �*;�w�k���9&Q&D�(n�Tk��x<
^@Sp8W|Y�*��$��m!0]�G�r��lS�����	����/mPE[��	��U�Z�Q�b���VO��c�Bhs�+?&�b�z{BI��a��� ^����V�${}5d��LW�c�ާ_A���D>c�T͍�m*��<��b�����.�hI��2Ϯ.���e�-gn�~�[l�ձ��޳�2�W���f!�o�kO� h�j�+��S�{]�l�ӈ�l4yS��6$����Da�Ɩ�'��9��n�&K6q������q6?62�0�y�����[�MU���n���a�"��Q�il��<���a�ī�L�%�?�ً_,�����Y�t1�������"	8r���Em���?Mc��@�0r.p/ƺ�
M�R`�4F�]=9s���I����rJU�s��p���$qcz
Ȍ�T��t�8�����e�28@<�F��������װ�<2�ă�����ihJ�>��ӥ$��?�<����9�����W�n�߹Rg;3�nz	8���'f���^Mu��H��E�O���.\k�Ç�a��A�+����׵��1^�@	#R����+�%HFzl��x�t���e�T���A���$d߱����*�J��^�%f2G}d8&���РJ�	��;+������m����f�U9/�A�BcF-��PC�3���C,oc��~w��N��/ ���Km��X�����A�`��������KZ�Yl�����8��HhIh���Ķ����q�ʽl�ҷ~��|�*]@"�# fEn���R4��%��d���|aw��:nK�L��G8I��0=��ќ�{Ҵ��B2��2�8�A��F��0����Sު��>������ג-7i�r��뫵LT�9�PyX{F`������LM�LTX��7}w�0��y��E�U�������Y����ً�XW�ٖR`h^�¿���0�S��w3���d��J \��,���X�)��1D�t�@螃��Ej>�}��n��^Ck��b�f�1��+<BcNY����a���31�ɦ�(���OI�r���L���`w�T�L��P�
�� ���32��B�7�z�pt4��'�> ���_�<i�mKX�G���¦�l�2��)Ź}�N�u�x����mမ|�v�j��sFX��r��ў�S�V��g^E�"��`|��+������f������e����ݴl��^����O-H W��W�sT+h
!6y��u��I2"��'y��ZH��_��<�q��`ʾ��)w^�!�m?S�Ģ��*'SS�ݡ�����El1�ـ��6(p��~��{a��Ǟz��P�Y�����8�6�!��U�
�^qO����ы���n��#%�My���� m����J��N>�(%&_���z�w��c���zx%��CnI��5Y�����0Q�k?�Â���I���P�)��1
�@l���4�a��}pb�l�&[%E7k��)NkL������^qNC��ҜRs��n�����G�VӴ�HY�a�+��VҠ
g��c�:�P��l�J<P9�����k�ru����qYҹ=�y4��h a�G���/A��tYI6��SK(o�'LUZ���7$�|��c�f�����ce"Mb�Q�뻗=g��<@M�i�*T����$C�^���0gb�:��1J k�,a�;+S��V�i������4@:C��8��>��.�����EP~��Z�
:Q�D�V��pwd�]�Mފ����֧nh�ǣG|��,��p1V�Ϡ'F��)7a�vz?J"a�ڏg8���V�'��[2��U��ϵ���w�����R-mߩ��4�[Hw�
���u����R	u�>�c����U]���9�"���g�MZ/:w����i���r,L������P4����6^���2�6уJE2��~��6�Y�p��%�s��|��W;ȍ���KbmF.#�v�t6����i�J�m��d(�\�bW��S����y�T��W=Ȝ�Odo��S�v��ޗ�t���Xq�8��� /V�mk]\��!GW���_�ؙ�O޸��RUۄk|/��b�Tכ�V�/>x�hHL�D��DIH�� V:��P�t@!��_\B��&O'�qCYw���ҫ{�:��?���`K��
8!��H�m����7D��n�
�� �<�v*d>�`����3�m���|�zD!�N�۾��9��r��k�!dqD�X��	S��a����,R� ʸ� SZ����Cڳi���@�7���*a6b�S�f��8����R���֕�yt?GTZ4����3c�)�ʄL*�_�dBx�gX�+�E؂�����6�T�x�q譩A�AE�%�^8�taڜµUB�OE����L�EN������H��/brJX�[[ؕ+>��q�����i ���D
��;5y�u�:1�nab�r�����P��o`��(�|�WY�S����4$�-�o�cz�_��_x,��ET�|�C!D��tMc
��*mː��'z�(���a���1u��ϲ7̴)u�x_��}w -9g2KݪLA�1w �>g�_w��	����D3���n�t�}U@�Hl�dx� �������bB��􈸟�lz�tj�g��!��.�����9�3��)�c�V�08`�|R��Ib�F�����t�������p>��K������Ըt��RrD�v@�eC��a��S�i4���E�˸����/5Pb�j��}d�N��5?�-.�������i����gP?��H�1p���X�PO��]��A,����A4�k��9�q"�/2fZ�ub�O���ɜg�2|S�įYm��f�&��k�t�BX��S7.
��utMD�q��7�BRp{����f
g.�-�RS�'�*�B�m��O����C6���3D(�	t�I��`la�������Pa?U?�}P�H�����{6��c|0G�\{�(÷zC�����@f�Ъ�_L1��8��Z;(���B�?J<�T����d�gg���/�m%"v8��G��{R�%/�nD�����VJ���^�{�����c���c�+n9��&��c+�0kۿ8�b�Ϳ��Z	$:?�^���0��ۑ�W=(�!ʶX`3��>EZ�u�mg����8ٖ6a{n���L,"�(�n{aT��,�����*k��u�Ƨd2{�w3X�FQ�E�T&k�S!� ��qR�]�4�c=�R�����mG�Α�`����oB*�-}GoJ�;�TI*��-qoB�4 �x����EUaC�����籲AU��.�]hgGh�M��^o3N8�}Ő���0if��1R�s׾fBY�+�@���+]gBv�\�&�]�	<�X9ͯV K�];���9��������Hu+�����v����2��`+&��t��/\9\���K���@j_
��an,�P������pU��ṉ�(�����&�A-�[�pq
�-��E��3kD���)9�Ƒh�S��Y��'�f�97��SA�?k�g(I��a
Ȕ������ٖΔ��ՔŏQ�Z�۳U���$���u�u�G���*�*��i#_�b�{@��������:�!
�HPM�����y�A���b�Ӱ&�$�� *���?l��#\���p�6���ө��ih�fBik��m�p�2	+7�+��R��{cߐ'"��+#�p�>i��`��C��B����ǰ�l9�qʟ�1M�\�b�,����z+��S�;l�P�o�M�o�����jD���ƫ���|�c޷�]���uwm�
b��2��p��dbF����d�c��p�;�\#mf����� :�<�>f��$g}U�Z�z	V������:�]e�_��ѼSd���ʧ����yG"�3�z�&]?#�v7�qӵ.����Ա��r�$��*@�$l�-�A��uCnN��Q�Q��p:pc�˼���B��%#���M����u�;&OGy':�9I�ރ�岖����AC�o`g��2� $©�i܀�	� ߊߨÆ�L<4�@�ױ�zr��muL}�;B;�6�%qU�
�-d�P����g��܎���j��=�g4��,�r���M7��Є����,f���s��H�Y�)����:���Z���S<a`3# dn���]<�,%o��{�wr�{�(�epZ�UCX�jJ�[� I���s�4�kOd��"@�Fgn��It�[�O0	hkM*���Hi'�ܞH��A-,JZۉ�G>f�y���H��
�`Bx>�6���g�[���)����ĥȗ�{��;����*��<Z�-4�@v)���f�}��0�+u�.�K�[e�,#��{N+gvd��vng Y��d���)'��%��?�:J@T��ǿ��'���}���I��׹D�	`��`m�5�1��:]��J�� {��դZ`ٱ�^jr0j�zLl�.o�0kN��&�	�.��&�91	[ Ꚑ�Q#[�����~3W�L�W���}��0f�����X\ �/��i�(�#)�2�������$�G���³���me�� {��VHʇ���Gf/�?pH�ԣ�i/኎�g��2̇9ZH�;�u:F�8"�Y�J~� )��� ����+�EPN�`�]�Jba<�J�?*�D�������!m�wUچ�/)�y�^OlQ[Ud%���Ltg�h��ga����#V��RAm�i������`B^
-��.\��s��x�9�$_kщO�']|����=��LF�6d��w0�+�N�
허^f�,�Ȓ�Tbv0k���1N���)ΠSUV?)-��W�ců!G��qX�)H�Ha�u��+�+�MJ��x���c�2E�5��ip�(R�#���dq�@�(tNR�_>�!<�7�Vv>5j�I=�f��+7v7�ߺM6ڍ�j�X+��ݢ3���#�Ky@�X��2�k��+h������"�ِx�X���B=��Ġ��\�y��>�^�ZJJ�2G��q5;�|5n�Ʋ�@�ی��(e¶�z���l�0�aC3�Ŷ��,O�W���I�G=_��Z�x+2=}��E�Oz�G�!�|=3�8�Q�K?�wn_`A��R4�D�*!�(�S��>;����~{p�{u�=wޏxk^�<<0��j-9a�G�p�$�Cp˭@��v���w�-a(	4���ޝ-oe�u*�*�̋s5��Ez |!G���m�Ќ~��c�� Ll��wD��sTd�άd�@&E1d[�Hq���;���/x�U �u
1�`v�̔3Y�_t��ƕ�(����������T�ʔ}w;�j1���L}���i6���:�-�E�>��{��b0�qj�] �8[?�a������������'9\�������R��@��{ż�Ȟ~T�i.�D�:43�rj4$뇄��ĩ���U�v�B��ͰB%ǔmB�n�ze}��6��[]�8vZ���_N��GO��,�IAM� ��WQ`=(?���ޓ��9n����з�;S��A����<xMV6�b+s7��鼝ưx����H�y��P�B���K�h�2�-/�h���l���$C!`�����#|>���֧��FE�p�7ܣ���g$�q�_4(�[E���O%Lײ}V��;��{�䳿�ܤC(�$A���n)��=L���˶�Y6�LAv�t�`�ב(��2O��;�������7%� ^�XڅYEj��A����n6ג�����j�L����|�4�է�ȓu�u޼a[/a;=,��q��%�x�w�N�vWR")BIj�����y�
���!�� {�`���t� 	�T��=,2G|��`�A�8�)j՝=�1����b���YDZ��mE��A���, 	b0��]��u���P�.� ��Cl��Y�ӜD-wߐ�߳���s�!����Ί�l��]F��� �o �O��؀�A�X�loF����qj~+)*B�Ӵ�Gjj�8 ~�� �ː�26�n�/j]�<�Wwk,W��M۲�Y��1;Tqy�9�1D�p<�L"�\���=�M����JHe� �Z jLǼ��r(=��3^r������1��I��@v��K�?��B��@4:�S�r�_��xi�ℳ���0i^)#N�|��\(B]����,e���"��|�k*W������Ŝ�2���X�����Kf�N,lSe[��l[�ى�@{A�Nm���4��$�1Q��j�w r� ��e���.h����|��ng�4�B�l����[{�ò���ɏ��޼،��j��<�_�J��kYiS�;|�p�2T����愁�p�\��(�r _�&:8�v���/'@V'Bf���i�$YP?ܲP�B���S�������������p��%��W�9���@�	��y�e�ű��ɝ۽��W'�|�#�؋(�?�JK+S����'�;�s�u��(IՋ��7���}��6nD�-�:�0Mwl��LITt�"��(Q��&P-�a"�O� � �I੩!5&���|A�:]Ċm��&����R�cYv�ѫM�j�8���)
��p,u�I���"���~LI��7��� U�K��cF��p�l襋`��=Ȳԩ��"�Rp͏Ѣ>r�ـ>N�������tu����>\N��a�t�3>����!4Rix�R">���ջ[��G��5�1�>��h܍+R^����BW�� #\�s �8�n2W�=�}�:������mhM��i� 3��c%u��U����>�q��bHv'�PPy��a�f���h���Z�=;�!�xw��[�}D$���Է�:!����P�< ^I�ٍG��s4���<{�'�	�����h���˰m0���pR�>��t�*�GE��J�u*=
�og��iFٯ�가�eB�.���3�?Фʛ(]^	F�[�Jt9����
�ntp$��!�4Cl�P%>������;� ���\�` G�k�=-h��c��5��V^;-ʮ�9ƛ2F����:�_��:\��3��#��v��#b��2�_-�	(5����5K`3�{s�_��3U9&��H��(���?��=��}���,�Pϖ��6��AE�6�C�� e��$=s����`ᶆ��\��5���#/qT�OXmQn	�n�z~���=���8[��B����Ml�� �T��"&갨�dcD���"���s�T�ۦm�^�	�H�H�����d�/�V5'y������H*��c����:\g6-�H�,]CEm�3�--�h�d�S,q;� v=�,%�ݷ�~:��} �|�������p���i|�]�V���5�m��2J[�M��
ۂu��X&nm��>��#�:�x�ɿR�s5µ�@
�f}1��}3�@�	m�Ub��i�j�V�!��_o2�@���߼�1����͂8
.�{.?���>�~vU��ގ��q_�M�9#(Wl�RJ�AF̉��v��ZP"��k���Hst�soٹ����fC/���#W>x��6�$T(���[ldD��w�VI�Eզ+<A^<��
H]$�7���wi���;���"�aD������[�|�;N"�N���8P�|��f�g�H���-/�l��7�}Pk6k��Tpw6T��f�' � ���~-�`��£2×�u^P�Ds�������x��D:u�����������Qs�5b��uF�t����Zy}Ɇ%w�ַ��M��M+��UW{�2��!C� �=0���<mJ�C��X�n���Kl:ZP�^ݥ�ȏ"ym���:����1�d����`�s0X�V�j	��?H�>��Ķ��t�C=��Fj-i�A��\�5[G,�R�����U�j�NF�y�+O�	^4�q�7`��G�{�k���)��+1�+��-&���iT��(���tlTh���]��A���~�[�m��o=	|^��ȷ%pC���h;r�r�4������Z��5*�ҹV����SÌ���N7�L�[�/a�3Ya����rX3�z�b���5lJ��V�:�y��)������IR������ջ����`�3E?�FfeLx�X��pD�Y�/��#]���B�V����c�'��g�J������}+ən�ǹ.r�+��p�lt<~�.eD^�lS݃-���CStF歷f�{g����H�R���S!��9V*4�	.\b����F��!b,�u@�����H��O�W���F��PoMY�|]��Bf�&��TEs�I�B�v}V-$��4�Oԍ�<?���U�F�L��ѣ�F�mr�����<�h��mN�H�N����Bg�3�A�����u�^��N��y��pfWS�=�QJ�?w�DB����˥�=�<�X�V�����~�d0\�~A�g��E6�b4D�yܣOo��I�qa�i��u�g�2H��|���8����>�_��_]?��c+�o��iޢ>����> �5[��]��wMw�m�f�I�{jEZ�o ���T�z�S�Zg���Tg4]r�s�b���d[Ơ���xG�`���%���i3'{�����K���g�=�Jf	�r8�>���@V��XVĚ�`�=.�� Z��jl��|�GF�U������RZ����s.l?bL�%1v���é�GFُeɟk��ޢ2k֞g�&�� ��qkqy1*մ��u+*�"��� 4��]���Q��s��F�t�4אtE��$C�e��p���bZWE�J�tcbg�{��.Ɛs1�8"j�|�e{UB.�ϫ.���'�m�k��
�O��-jE�	�ܩ�Rmvɭ��1�6d=K�]]�~��O��=���9��َ���՟S.�U#ȭ*~��g�i���Y/
3^N�m%�^����,��Rm�Z{�bV=�0�1)?~ğ���a U�G��q����u�Бt�cٛK��t�q0�,������L����i�ZM��YO�%]	�A�)�v�|���RD<�Z����C-]�7��|CX��4/K$|�Un&��(?h�������N�J����l��੫�Kh\U��]a�6�O�����#�����RX������lg� ��:�HN?K"l�;���{n%�s�����'D�0!
���Ԟ�~SdR0��9�'�?%�\�[�1Y,���c8��O��fM7v��͝��v߾U��0[� X���<����d������_H�D�0:�}S��B0��ꀋw��VZbk�ƙ�sWsU�j��F�T)=�H;���� �9SKKߓ��4mmE�GI�c^�C���w,���2�і�����5�jMb�H��R0��$tj��ν�5Gc*��o�"
�>	�p�,7"������}]iV�4hZip@�p��V4>(K7ځ�8���Vq��Nq`���uD{*3�D����m�GF��KCl2.�0��G�q�����}��La0�c:�P�Tv�y��Täh�b@j�o>�J��Mι���u��O9ƽ����^x�}9�]v��E�'�m��x5W�O��R[T�2�e�����C5�zb�l���Z\���DW�ʗ�f���-��������+�(ު3�>�$A�+@�/�<PgT�,����U�i���fS�WAs��u���R���P�F��;ֳk�R�ӏȉ��0���Ͽ˿#����L
m�F"2E",�*���׭�fv_��Y�zͼ*�$�V��-�œX�+��)u)%�+yL���H��W�PJzb��"T+w|���]<��g}��U�&O`�o�w	�
�+]�=��Xz�aG�G�X��F����,p�� ��9^�UΩ���>_*����*��S"c�K��׀��	I`S������T�b2�Ѽq<����r(�˜��	���?�B�Ě�����>>پ{��/o�M(F?屻�]2JO�]�#��=ߞ�ų݈C�h��Gj����+kM�L��>�H1����/W�N^Y�dQ��l�W~e��G'D�2>0�uD��$��ZSd�kd����K�E.�~ۑ�.G/%5%��.+�JZ�SA�����0���A���`-���.�L�"�0��(Z�PJ��^T�m[W��	�׆��B��w�K�l�Z0д���Lp�Y d�9��i���KA*ێ�XB��ތ��W�|��.��\*��r�kf�-Q��b��=jj��߿�6}ZY��$�g���om��5H��0���ۼ%gYE�C��D�\�-S�әgwe�(X	����i�+\U������ɯrVY�93e���N�V)O{�����Z���x|���%�,Ȓ�S?�.j`���q�l�eօo�/���n"k�jݛ�'a�t�*��,����H��=�ԤU�l_�KW��+��d�l��2���I�;�	�Q��Y���f�¸=_�i���F��VQjX=C��>5���4T�ư��;ĥ~����G��5S`�椖��K���f'��`��*�A����E���i�l� #��������F��0A�I9g��$��Ը��%T�7���|^�%$�%���ȁ��9���0�������V���Т���c�m|O�@r�&MdN��i��Jջ�{S}mK������եA�Es�������w��)�sbHs�F�a@������2[�0��� ����L�b�I?�32|O�[X#1؃�~��[�D�ٗ�D-aZ3r$��юc�ً�eW��+���l�?��g��\�IA�ޖ�m=���ô
�Ed!
�{�9�����ݒ�w<�R�>Gj�̯�^�X�?�nG�1D���*�*���-�����n��[�[�1n���m[G{Q�oKx�N�T����dhN�e�[�̪ A��;�84x�{��hA��+�F(Нr���b�d��߇�S����N�/Oĝ��_@^�>R?8Ѕ�P�KHWa��w�|ZX���I�H�d���FJ=���F�&a}��c���h蘕�˪��e�q���Hv=��q�����S�'�ĮX@�f���Hª��a�1�i���ӊ�??��F���g��{�=���E�	$��Y��/��/)�iq��a��CFO�e5�l�E���&�}�0���D���O4+����46�U'l2n�����\�p�9{A��B팸1M=�oԚKL���ꃾ�m�s�f�j�IZ�u�#o�3��3Lu�p�%�ͨǻ^ΞӠ,���yj��_"5���D�P���puԤ崁\�T��B�9#���S+5���YȰUl�������U��q�[I�r�sV<��c���[��ʎ�q�}�P��� I�����LP�=�8�Zs/"��98)f��7�j��;�z��^d����h��Smܰ�Fb������W���+�g��2Vd�LL'��p�0x��`�3�y����\����w���2:��?��@�ciP �w�֎Ӗx\,���H����"�3C=uΨʠ�R�h��:�v�cBA�k("��o�p�Aҥ�iә? �A9Ӹ͖q�6|���{��Aӣc�L-G���s>���k�R)�A;/ȃ�i&qx�e�!e��=#�Tq2`.DC��a]ȉ�i�9�R�%�ê� �:��y��˞�Z��U�9�KS��Vy8gp'
>&C��-N1׌ձ�h&֠i���B��U�b�m��|SW;>�^���@>p�@�NזXz ��s���鴚����fv�C2{.��r���0�d���0�Ɓ���6�NAo��v�S�(����,���u�v�0J�Ɗ��N1�B� �1ܗ�t�@oF��:ۜ=2L�+�G���Li�9`I[��KN�r�U�(��3�b;^%߄ǐkh�+m�����D�{�2��>j�c����sԔ�vV�Γ�q�bk):4?��@~r��L�TNx��g�(��f��ꡍ�8���o(i\��H|�]��7�� a����p�f��YD��Ź�Z��4���0�,"��;J�2h�U0 �D5���FW��2����7_�Ɓߟ�A�oޙ���aE��_Ǵ9�����f��ɑs�Y�נ�6h�(N��H��x����y�n�G�����z����ǿ�3�����V�H�/�D���|�k�1�+Ȑu#h�-#�(�/yu�6�����c��Q�P��?�Ϯ�E�J��&�@Sه�{:�$m�tc��e�9�"�O�yjHK�/t#c*�E#饱�zX�~��Ň�"A��t��><�z���tx�Q�����qq����p��Ly�����+��sw��[����iD?�m�X�4��y�;)�c(�)۱����}^�U��hM�`�fU�V'���zǒ��x�Sy SHk�������h��uͣ�1�7�|3�Qk��łbh-�>Ա�4P�'$�a�!�F��W>Ћ"�M<������r��T=QMѠzJ4qsD���s�	�*n$��g �ȣ�E|'8)���̮��3����w�ޚT��P{I��>��}���ȩd������m�����2�Kg,j���7�ߟů��yi��#�H-̆�V%�9��Y˸����E%�����|}����]Ic߬�%2���o؁I=.}h��ysT�V/�,�V=��� )�����(&��違�Zv�4����ܵV�@eI3{�����ɠ_���3A�z�Ug�Vr�V8���$�Ak0pq�bQQaip��6�?�Ց�%�QU%�������:�BDa�$��8h�&�_ xg����ҟVq���9�QZUj0������F�:�P���][^Q��c���)HT�uO�������9�v�j$K,��=<�(2�Gn���Wõ��H�<p�k�5�F=����yÞ�#}hA�֧
b�����>��=��-�ɪ#��L�ldu:�zS\�F`(X_h�=�3����>���$9欜ݷͅ��e��.e�eUjxt�ka<q��{4�< �Rgpoq�D[l����a�{��0��Ti��M�f��5W̅��&��HY��������O�#�����P��&���q�К�-'-��QP��� X���+yVϘ߆�2C�ޘ�R�-�{���UY;&A�6��Y��͞56�������`m�%?rB (�2?2�<��B�0s���d�zNJZ%|L�Hx�����Q�ӛ��,��wj8�(4'T��AT�TV��+!�+��j&!�<J�Zm�ÿ��� ��:�Z�m̓ԽZ��P����w�X�d�$�Yt�v�U�7]��T�ʹx������` �P���*��{Og[�˝P ���m�z'�:�CL��	�x&UT�'�p�����}޲}Am�f������y�G�|��^��C+�)r�w��K����e�c%����nG@(C �UB��8�^���X�]P��F~�-h:�"r��>�0��M��-�E����Rlgat���<;|h��;�H����-x������RE�t���hC`�n�\�,|a��Yy���!1�����Ⰵ�D}���G�U��{�& ����,x� �Н�9M �>j�������u�)��|X��L�׋7���O��9[ٴ���#*aLb�;*N���sa%0���&�,� �t��K�+��*5c}�v�N��$��S?��ó3���s���h;�r�.�Y�/.`��GF=�d��U��¶�E��#����y�c�A��fu�~�Q)!�>@v�m�{I�yS~=#d�3�u>le���p��N��_���oI�R��~�Ɏp����bD������7�c�*�i ]tsL�������c��`tϫ8�
=�2���^��K����>Y�s��}����|@��u~�y�?�6C�Vr}t^��i��\p|0�~���u.���
��M��h֪��x;�����	Je`�x��> |�$��e��oq
�8� �Y����]%��	��.��&�`,��W��`��͌oȱ��9Ϧziyg�{mQ`��o�o���rbv���N��Z�ѽC�2�]U��4�)�F�����YWm� ���_�s���py��r��0C�) ��~�w���B�m�T�'"&4��G�Հ:f ᳽lΕN�,'Tj˹��ͦ������7�S��2��X�!O���Ի�
;�(�}�����<�s���]S����'�����؀�{M�|"T�]26�)�wvd���e;�w+�����8+\0n'clz�z�o^k��7`Ր*�S"��,s�.�1��ߘO����Zb'�&
!J��?Y>�T�TB��R��=�+��I� �$U$^/�h�����Ɂe&*�/By��"N����j^�&|��&T���\��t�=4��zg4���VY܁F�<�7�h�Ʌ�a}���z��9�66�܃U<�w��F���$�}���FfZ�*y���M���_�_jd���|R_����\�JZ�[�jԞ�y�ig4�|����k�Hh3|B
�$C,����wO�c@��qGՐE���8�f�����Y�꼾��-\�C�U#[����P�X1�.}������{�n'/.e��ΈM?񵥙^>�a���@XX����.����4�щ����S�a���H%!�ma���(u}��܍�ŗQ�Pi�S�a�Ǿt �=7*
X����H����ߞ0 ��u�°�(�Kg��� (gN�����nQ_ ��o��q�0�W�t�I������ ߺd����n�ed�� ��G��HP�m!!��q2)ET��u*�pY6��2�p~���,��s����#wk���y��O9�pl�R��aY�,��m,-�O�!=���j�d-�-�O��	�}� M�T��'`qN=�t��(�ov�����h��$�5T��V���k��ak[<p�bsA����	���Ѥ{�� ^�h���ݰ�-VR$\��y��eHC��:<�;JrMl'��1�ǡȩm�پ�#p ���)"�PX �����oo�`Oo�C��B����wT�v������T�od��׽ЪG�������9*� r��o��C�R�P�-�4��so�1�d���Wob��V�K����H��C³Qt=���;=ݧ���%f�s�V�B���E�-�>_��o�-ۑ�A�v�{.���G&t�ޮ���o�1�?�-��s�Z��v���A��BA��#7bģ1腆`vGy�6�b&�\%�|T�0-��bf8�.8{왎9����T�s���D���i91W��v�8���{�[ezN�������17���a�� ��f�,����+�j�E/�&"��j�����)"�Jf3y�z[�lKfHlsՃ/��+���G���(���a�Ʈ�9����slڈ:Z�kn�x���%o�[�aB�F�f0w.�*i��n�%r�Ґ1��#z�5i�"�[���H� 1q:��%��6��p�7�r��0��sO�Ȱl(��z���.�;�����H�t�����s� �N�v�J�I:'I҄�W�S'��d�r吓B���=Eq�]=g>hf���3��l۸�̣�7�.�*�ru����BTb\LBT�SNvZ*)�W��,���3�YTB9���3��'���D3���G(`�l����٭>q]̠�����+	0A�x)E7%�u���@ݩ'{��p����!i���e�"F�Ƭ��d]!,�_���_�7���F�dҰi;��2h��4��5�����ϙkQ/���I���h ���?8�݀�G��nƎ�])?�P��\��j�����b+k�z([���Em^��O��
��T疣T��]R���ɛ��K�!��f~�Zl��h���Xv8�G�ſ~wG�h�!���sEO�ɣ�C5a��<.8]��n6hD=�^:G�{CC,@����վ�J.��:w��L�'�ٻzc1�aPk��0 �ǆ�r��>�/�%��FxT(�=7�a�L���D�Ft�0��z�T:@����Ǹ���cy�'�̟)B�8�'�s9���]Nx�G���S�Z�3��T~
��I\�sC�q<�l��;�9�y��0�ݘ�^��*�����+i;�I��d:����	��4,A�2��PA��v[<�H���D ����9������;�u8A3����Yy�KC�*��z��sͼ�)����é��yI�!���	�p�D�����U��H\���yɷ�n:h9	)�-�WD��|!/x���P��.����B�}0��+u}��H�[��g)�ZF�~eB&��'�ڜe_�u�ۺ1�<�?^7?�h���H1L�w�������˅���I�����4�	�+._��;��R����X��$3WiJYDS!�j�M�i3if�uwu�r���p_&�yec%��}�﬷���"PƂ�0bf�L�[���hpD�Q�(���������xi��t%=�u�@�A}��Q
WҖ� N��=F CEX��I�b��k�I��5��N��c��\ۚ^}9L�m��Հ.Zb��dz�⤇Zx�ɋ�4�JsjL�Fo�|2͞ٺ�t��'n�g�)�ih@����rL�}��b���bA��}�&,����BFv#%�5:1�o�o�� �-�=��I:|�w^�X��X���+�M����<9��?��G=w!�"�U�>xE_�n�G���A�к;�@kk-�x�ǻټj#���1��������+CEњ`�ޫ�`�
�G�~�ڌ!f���i��RX���1����jb���T��U�*d��lQ��7=o����B���F��e�H�=~�f$5d&:���e�����@�J������p̼�|:��3�?�v`g�O]{.d���(��')�S�J��~k�ha��A����2�\��ǖe���P�B��``?�H����Q�jD������M*L��2�/�w��a�<H�|m�vY�٠��.��CA=����t�J;��<{�JP��_½����O)I�S��_$�wiv�@ބ���|��C)z�B�ݬ��)�#L����ޘ��Z��;�Fj��yH8���o�L��r�&���J�)�tJ�:�ΐ#�I���|"��/hY���nU��B����A�T��ă�CS��b������	� �!��.�a�@���ڊ"ہ���Ue�z�'��<jL��1y��"��Xu�h��=���U؉
��W�iTf�REB�؎�J�X���n�TgӵL�!�L���eӋ_�S���> �O�,���3|!nIhuyr����� hAs�n����[)fX�;2�MW%LR�}�r8<?i�f�P���T�� ��w�s��Hg�.�\���~k3n;��(�����ko�y�je���x���;�	f��\5�t{�hI�h)&�陾9��Op#B�b�Z�L�,���O( ���۹�i��_��D��F�t�mXf} �`8w�N$�r>�6x�#] ��9�4��}�kd�T��������HQ/gr=��Z-����7����ȴ,t��	���k���������<�d�n3Y˄�UX���āB0�8$"���q������(�l�f���Z.�7A_c)J;M0C��y��� � �x��=�T��;l	�a��^E�)� �-����n�y�8�T?�!RQ��Pp�*i`��S�7*N5d
�)&Y���_�U����A�ZH�}/@46?>���d�/�'��H� m�k=����t1��"�ᗼ �w����`�Jr��n�:j�:]ő���#��eܝU��P�U�����N9ww�F���=�;6���!r��|b���-�6;�x��!���|���[�� I�)U�C%�
�8t@�.Z���{w��ȡ��@bx��V�-]�k���kМC�+��U�|m���Z1�Pk���aL>�:�ip"��k�`{�5�7vL>O��M��ί3�!s�*�˔o�C`&D(e��qX��S�Y �Ӭ�j����Ղi��[���y���g�z�v��yE�sǖ���!}����B���U��k(��QP݂���~Io�35�ϐ�����(xӹ��c��;Oae h��c7�<��w�,���=⺸=)��(�w(�����3���L������>�/�H�Pˀ�zR��D��F�����骸aw�O/���H����[��$��z�L�nzP2&{|0�~�!�
_)1�d�B9���[��j\z��p^m;x�>���
 BHN�����إ3��^�lZ ��~���`��ϵ�EwLs/�"�gi�4�[��|�UpB���1�$�]����M��[O+;��hߏ�kX=}��7��Y�O�G��!��1 �ڣ���G4��Ԝ���|�QU2�k����z`w���j�|��9zm.dD�bDg�������j|䱋%A��?s��V4|?ȸ}I�����#����o�t�d��L��e��h�hw/-�`f�r���a)�?�i,�S7Qǂ���n׼����4��!_2w����֞>{G����O�I�ss��+��m�����(8���A�ս-�2�Y=au�q�A2n��ܻ3jн��ݜ�4Hfy1�90XL�\�E_�$w&5A��D��K"׾�}������I!���ӝG�+���.}���g��	}D���sa^��jr~%��X��B�*T��Ȏ	���#���G�TB��:j]��*���I�ƭ0��'����w���u�ص�8�u���(���,<9h�/��	��E�N~<"�?�ߩ.`�BF$��z�g���Bj:;�T�0�d91i>�Fh����J�W[,C���]zg6#�jQ4� ���qr��PU��µ;���i��M��>�.�cw�J�1��{�F�v}u�/W:~~*5����H�l����p��P/��������|\;��@2l�䭝������ތ,{�N$P�LA^Wz�#v�f�ŗi�3�V?�*s�3�0�?n��P~;T��`.�
�]�^5�9���1��AK�+��Y��VdGQw*�q��/)�.�-�����+6���Dh�K��D�:�;F�$7v�Cw�~���-�Bh+��r�Z��9������L�.c���!�#��X���P҇�
#(�Q����o�)P���&Db����>�;��^Y���x��6Ce�Ci��'� ə�I��y4����#�T{�� �Jj�T���/��*��C��jq��F��Q�=��wS��G2����%�7�:�k�Y���i��vѯcY!6���--��΅�TWr'Qܿ�y���#$h=g���]�9:��_������2k�߹��<&.�Q&�Y~h'N��x��k5��!�]��A&���&����r+�;N�I��E�g��WW��q��)��D���8}>��7j�.�MH�WC~JLo]���9:<���p�&�R��������$�lo�g죜sƄ��]F��y� 
�L8n����n��Օ��&G�b)�y;�l��u3�Ӧ�}�t$�	ǲ��/StX����.OX�JQK��UӤ�2^�RJ��6Hҋ����:��t	�f���4\�	W�k��h����f�$6h9r~���ے����ZG�Dg߅$���#Xx��?����PGV��K�.�����d-��S �-,�Y����L��hlt���t�T�͠����v���Q�W��~��Ǟ�2$��E�����t�b��g��L�x;��������ja��#����S��}��zy]��A+�6}'�3�,�/KE����B1�H$>e��+a��>-t��㻤��2��uԟp�L[�ݳ%�*�|%Ie��
`�|Pi���\�@n�)�l
�4UD6^����m��Tu��Uǐ�-5m>r;�Ma�rð��3z�;�9J��)��#;���7�R6�	��i���B qo\�]���t%e`AY],��G&���{b��=�ve�4��ٞ�Ug�|!/	]yK!�	s*���-D(e�{����vc�*�LK�T��H�h����g{���E���hIsC��WL���W�r���(<幓�dYW��?�6�ځ�6����+Z4w!H�kd�<w^�~�t����8JJ:In��+���m���j��h:e�F��a��8
S��ח�������������غ	�����]��l�����J�'�w�xX�G�:�~�)��х��̒�W�j��I��-i.�G��[$x�wuVH��t�s��P�\�;A�B$DA�2��#P�w���u٤V��E�o���*sVU75�I��Y���;��C�����t��骬�2=#/�Yr����kA���+�_q�>!A7s�Z�j*��l�'���f��9[囓�������%�9la����{v�y�������>u,$�Kg=������>�,3�˗l�+�e�&�Ub!�~��|X�ESȓ�����I)}�zq%g����噥�:����/�u6�ń��&1��MÒc�+�r`�r��g�����	/����3%���K�"fFb��Tl��뻙N�D�J�� jD��R6̧ċGJ��t���W@Gc�#|r�*�!Υ2Md��|U��z!4Q�W�_@�[�Dug�����Y^��l���̢���Ŷ+�5@>�H�C�C�[�KCH�o�3��HT�Zjz�o�vZ�9L�n'[K�`E�Wv$�#���F�h��4������'Ó� �Y�~W�%R�(-!:�D�wξGb�J��k��1�v��H�a�u�~��+!1)�^��G���[��MH%l��vG?0��ā>[�9���&c�Q��P�u�Gw�C�A��U&?ϖM��2	q����n��:��������hTL��@"I�`R�3T`"��U_�o��^0݂����Ly�umZ-�M��OkT����	�"Ɵ���  -5��z���侤�7�j�{��|� �mMZE�jIg��,��LVj}�OU���+/�mh򥝅GWw$	S��?h��{��y!� G�����5��(�rfrhfi��8���P0l��;�#���u��'5�2�s/�}���?�΁(l�R��^��ӷ��UQ�	=��"�/Fy�|���ǘ��Y��l��e��ű��hKnb�oTYGY/�Cu�'�@�O*���QD|������M�Xӄ�k���
�����~_���aD��@��^���s$i�8�3~MfQ��^]����*���m	-�B���2
〈��1P��[>.�@�=���z�c�{��3/V�g"�S]�M�z �Tn�����.�a�ϟ.��;k��՟�7j �H����QokТ!���b���Lp�U���������)�˫)N �)�p�gKQ�	�dby�)���Q�������`�
��~�;Jڕ����N�;��|D��^l��r��oJƾlސd�gM�d1���K-\���}w�8��[[�7����s���塒�TPb�&mb[qar�#�j%?d� )�{��#�/����K֣��q�����1ZS�<�Q꥽"9`�=eW�hzu��~�,�D��o9%`t��.�8ƳV�b��̓�.���ƼV�6� �����t��ަ�#I��+�^����B�D���K� ����ަ���׳�:�y��7�z���A�<� JS�>���{�Ԝvw�{&y�^]BV�c����5
��+]<�m	˙Z�_�����Z�.d�=R}u��g���ȳ�v��r`�*Sc>j��>.�WN$R(��YtL�!j��a��c���a�Be��_�u;��g��@W n?ɩ�Cb$M�~6U݌�XD�M.���1C;YH���i���ܝq?�%U㮚|����.�����Q*֝����u�V����oW�����t�[������N!�.1�~��I���-�KC|�"�YB��B��1�vSm�����!����uM^=UgJU�ަWI�)�T6k��|f��ݚ�e+�*��#�=�j���}��N��?��ǡ���WK��;�~3�\���кo��N9�0����w4�o�w"=�'$Ç ��K���\3�	���ĺ��N�[�}:������	�3��_�?C�a��9��z���0I����`Hv:�\�^zA���$j6���������S���8�cc��_;k���TC�����_cSy���%�~�{?Jq���6� �ɐ�a������y���PSn�覽�Q�l��O��LZU�-]���N�ܡ��`O5���Z{g�˟���}P�Mc�:�p��Ș8�'x1\���m�������~���r?�!�J��IP�pO�ݎI�G�挑�pZh�������L�8]UΑ��?�\�6��(vP߫e��Ђ?rI0��@+����G�#AhO�hl�.�em_+�P�YWY�2u��O3��:s�Q!�E�����HCNC�⑈(^���3P8+
�a��`�&紞��um��1W����5o)f3ea	�A���VS�a��)��1H4����i*@��ݯ���e��0tjl��XI�[I��
$�{��d��.��M�@�[4 �i[��m��ֹ"8�Y�od#�æe9��O���	^�
�ʃ��;�2�W��xv�/���N�l4�?��޻�qn�(&�?����7M@Z����������m��;��	��T+�iJݕ�o�N�r'��� �8�����1e2S��\��$qv���0�pP��	� ��ǹ}��eڝ㵝S����ġ4̉���q\�-�
JD�6�iѺ`){���9��עM��(��R?�vO%��� �i�J�;x_y�Pǩ,/�a��K^Ƃ{u�����$�.{;�f!MG�X&�|�