��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@��D���F�Vp��t��<'T�z��o�ބz��{�s�C�Dp��-)DC��l���%X)�by1���:6�/+TV[��i�b墟]d�:��Oa�#mK7����ZT�+�`��Up�ZZ�wC<H3�ؔeN�r��<-�^��p����b!�7����t��lG�pـ�\R�����Ǚ�0<�r�D~�X{D@�x�uF�
�iY�5c&@�ک��
�#M���)�N�w����S<g?7-�@�ٕ�[��p����lx��Z�d-$d�-��Sp9 +��5Qa�<~�V���1F����� �4�)���2��&{<����: �`0Q��2.	��CX���w��CH5rP�D�<�r���{\��h���a�ө�YDƧXI[�d_�pWA�������]�k��n1��>ͥ���^=F�5&v��I���J@^D7͞�E�$V+O��=�}���xܠڦ�E�����j#�q�|�'��)HJdV��R�_f[sWgL�����y)�"5�ۜC�{fᵍF��11$��g{Oc�&�"�]���
��A�k�S>MR���܅T3A%4�lO�L��.��_��Ɏ9��;ϙ����g�h�v�RipTIB��|`�\��q��0�!�Qײf�2f)ְ`~S��1~G����E�aW׼�4������k�*Q�~צ~��E}]��t���*x��_���4�*_z��-��ǕoP�}z����VFʶ����T� d�CP��5�D�me] v0�U���_�6Nh�%��3Y
������J=���=�#c����0<tZ�ܫ;\ׯ�k/�tJ_�#BJ=�͵U�g����G ��"եT������6aa���6O���8ǉ�:���$�ۯ@͍_���S/��e�{ϼ��A�A����q�!~��0�ɑ���F�7f%�B��������yJ~v��=4/�����CP%m��>r�����`M(�D,۞Dcc��h9�i터6�}����?_eV�JSc���5���**\����A��?�EJ=���ƆvffFT�2Dt!�4u�]BC������;�de��%��	a�9���+h dn�f��`�In�R���-uc�(H �R�.SL-�^��꧄��$d�m���<4��b/�I��[قf+�	?8�nѓ�����	�z_��K1��(}��%��dò�1�NH�B+X��x���q�@�(B�z��u��2~��(������n�*��Hc�e�ښ�_fc4۽����2cG��ڒ����ظ6�c���^=b!�ּ���e:贜[m�5� {i�"�?P~VhG��Y��R�۩�"��Y��,	@A�+�+��	���v-	���hR��}�����|�zl��6�u�s�u3�e��ƞ�	s"���Y��Zly?�����|=V�����g��5#���ǘ�,7���8�vP�Ƌ)+o4p(W@L �i������i�6�r��Tc�П��GT�<Mk��V|��Gs�x�5�!(��ux���`1bO����s���$�^{�'ڟ��4���4��pW����iic8��m�?�$J7�H6����[�wC=O��������|�H�Q�}��f�84����G������I�4�tʊD�K����B����L{]�h��9�*��4
9���TA��J_��7���t�q��|�O�n*�����(@�$�G{*�� �J�^%�{ʡMU��]�t"��Sٶ�WJ��66�^LlkG�K4%b
d�s�=TkZd�Mc_�q%;0���&��B=�#����_���'�ҩ�7��.���/��̙Va��5���C{�/��7���D��(3j���ԥ3?d0V������?���T���Hw��!��c74:2_��6
�h�^lU$�q����P&�I�� p�ʴD�KX��-r��XRP��.s�N ,YYȺ�ኍ��O)γ�oF�E��l��ɸRO}����rfq��K�v��#Vj�I����/a���՟�bN��H��j0����{����l9�='��+ۿپ)�"|P%�(;���Gq�kR�!6O��eF��sI\����R}�B(
�'O�_�E]���c�K��U$/T<�)|��^u�8j�+��kA���g*^�o�II�{��f����v�2푰��=Au��+͔���6�)_����4�&�Cv��O��ݹ�	��T���2���@��Q��Ao1��mS���CsӇợM1�)��q;�OLK(��$�P���߉;S4q�c͕��X�B�i׎�Iф�b�Vic�X,Ĉ�S������M��������6=�pqp"s�S���V8�b&\�j��)@�G+wQ} i������n���]1=��?w#H���XiҰױ����
��S̙���@iqm?o9R�M ;�|M�-���I�!�<�C���iz�ZQS"�"�y�2\����^-����~#L�(��Jac%��*X1���s�@ �?> 
4})��:�N���p������'���Ed��GJ%��׶��<��_���p
���bǆd�
��U6K���gz!���wS�zo#�Hj��y.Iu�4>��8(e��>B��A�'`ܻFY6�vj/�����J<rR�Yk��PD��5�q��ŀ·�,<�P@MOT\t��ƭ�����3�1����+�����N�'_�IԺі<K/软E��꩜������9���{��0��OJ�f;�(h1A�&���H�0�B��n�R7��v����a�_�ޗ@�e����_Ӭ�^���#<��]8��*햕`
�˥ָ
��Q�ⒷRA>���Iu|���C�S�;5f�7��8K7�GGXåƶI������w���+~n��#�� �7��8�iu�����^&�e'��ɨ*����5�4������B���:���xc/������=�7H',����:ѥ?�8W{���1���w�0N�V&���4��)���u
)+�@�H�y�UP��v�,�^Dl=q�m��uiQ�K���].B,[=��Ԛno�����0XZ���` 8ba-O� �� �ôS]Ȋ��0�#��A^�o�},?��.��i*Gw@wD�`7��#�����pݥ0;:��H���W}$Ǹ$w 2oD����v�i������]�K;�������������]�a۰֋Q_a�v��D1o��6��T"�����厣_�|�@[L.�dE��O�tCd�S1�{&��C|N�O��	�2z�hn������ೝ��x'�4C]�b�{��I��\��(��Ղ�hE�"q��M ~ �,!���%n�! �Y�{�9�oY�I.��-��V�����]L��E��U3+���5���I���#?��I0���)���D�������/���B��x�6 WV��S���{Y�b����Y8��i�bcϐ!���X����J?OӢ�pڳ����=�9�F?y�3 Ӌ�[�l�k�����R>5iw���a8��h�ΉM��c�"���2A�58>�ru"��$���Ҧ駉}׀ҤH��Y<���ǭ�a��@D�PF`I_�v��*�[*� ��^��f�-
�����H=oB֫�?����[s9Fݢ��})]�(�^t^P�&跊�v�������q�]�<��uk����+N��ؕE������ۧ��'j�^����0p����2�VY%|�j8^���uؗ'Ԭ��=��� Ô�-��S������.Yي_�Ҹ�	�WI\����U��,��of�#127��R{�|�2&��|�p��*��#����5��A�������=���e7W���moh�PW���x�r瑚*kfl�%>�6��Ԩl��h�>���CP"Rf)J���b(��3aab�u�G�6����v��o�l0m#e�@ZKI��`U1f��ޮ©��Z�"���~)��V}��o<�Ez�2��`=����dhAt6]�-8�4��	O��RǁR6�5h�;��,BM��ݐ�.t�����q�7WC��1 �SE�A�]�E�n���H�V/�F~�6���s�����-�^z�cQvJ����}7tw�� +�,xY5�p!#�=���Mտ��na�c�j�MavR������IMf��Y������=Ӻ^���E�CVA�������_*�,���'��Q��۳�b?�3����on���k�h�
��G؊�ӚV���crgY�ս�2�iԁ�}�,�)���8�x�#ר��;nx�+�
m�~�N=���دj��r_��C����(�뮫�\��f��w�&��3�]M�S�@%`���L��:���6���M[NBi��"���+��ԷL��������WU��������b*�P�#п4��-��4w��:y�LZ�Y�!�#Pt�AZ��h�ꏥ`VW���.$[�m��瀠A�S�z��.��j���\��E1-�9�"ʇ7��U�����B���ek��d	��qb�aS��tӜ�ܚ�Ո�G!�3�S(�����3!-BE�M�������s �᯦V�͏3���%.	&R{D�sNY��Ք�FJR���R;�aU@�|T�n���T_��vr;4�R�$��i� �u=u-)���<��g��}ɘ9�:j:�U������oZ�Gճ�Q���b!;N��F:��} ,B�^ H�<��5D��߮5@��������s�Xµ��mC�m��>�Np����5p��Ps�9��� �v��o����Bh���Y�N�ի�tޘR�hԵ6�1f��.4��0&���(v�ɧ_<j�7��e�F����k[�C�w(�b �q�B��,#�t.[::�����à�,_�(2j�1Ģ�<x4�,��U\9Q�����_N��=��A�=�K
����2!`8�ŭ�����@dU��b�bq�O�����)qH��y��&�`����Iv;��%D�P.���&�cT��,k$�ze�c�Xì�Y:���
�&�f���I��_����:W3{�Z���]驢Ac�b̿?���~�N�{��|w�_�ſ������ע�@E���M��}��d�p#����z�������@�W�R�;v�W_z<�a}3� 
�5�C��'l���׺M�C�r]��D)4�0��I�����I�D��x��0�a���d�+�"Jl��k,����^�_F�/�r)�x�"jf~.]��ҿ1����܍���ҋ]&ܛb� �o�<�b/���^��}v��	Rġ6��^ ��
�6iZ<�ߔ�#|Vey2�ޱ��(�f����w֐�{(�/���UBE<Kh��xX���ܐ��<9gk%���C\}�u�)�&��w�Ҳ� �Qk�vݒ(�$}��ĉ`���?�n��F��ȑ| ������˧��5��̀�(���� ��p�h����*�5��k6:�nx�'?�rY�d�h�A��UY�Kv��B�����"������/�	��$���$��غݥ���'��������*TXS�;�{�Fk��V��̙E���Rc6��d!Y�Pg�ߘ�:gD�к2��7�+	м{�g�u�P!��>������V��P	��(HCP�����}\x�eS�	ð$���rN���&V#,�S6�*9ߐ�y��)X��e����%�y��"�r�}Zf���Tp:���Խ�w��0�]��D x�|(zV�H|2\�ඛ⮱^὾G�[�`�)ё+������M7�,/�ُ��պ�~���	Z��yk��C�=j��Z�ˋ����9R�^�I�^��t��3G�SI^m��vW�;�%+'0
��f��rk �����9M��X�I��TWb,� ��^z�����i���?�k4�үM8�\�� J:���1�X�IW$9�G��a#�)�9�!��2v�I᫇=�������U�L9}���ث}v�}�[�7�~[���e��$���1eqsq�i���M�%�Y��J&�c��P��aB�Y������:8<��=`��R�آs��Y6�Sd
azȱ������ cMʦǿ�/_��b��+c�,�������*+gΪ����&g�� z&�!S<<�]ҝ~�ޓF5.���/'B���G�}z�P��˙��i���j�vm� WL�U��ڙ��V�E�� � >XX
�G<�T��-W��v
���٠��F�Ss���b,,�߇�vφ� c1��t+\��3��� ��z�a�Ei$���H �8$�+R���;i�̨_��M�w������ul#:��"Uŭ�A������m'��V�i�6���Or)4�04EC��rP$�45�#�~���֛�J�-�P�F�'4�N��:������Q�u 6]�a�ͱ�^bوO��Z��ݹ��lAy�G�b<�uƀ�wwrd;�3��!����l��a����'������R1ǿ��8�#�#��+p��m���^rfd+��:
�K+���Zo{h-6%��u��"n�V�H��H��VZ�cw^ܶЋ�gj�z���8U����P�6�%J䥱������T��Ʈt����RI�P�@�����f����Ȭ��O6�}�H�$��u�pcZ�؅$
+Ƿ��v��ǵ�P��"܉�/��A���+k8���B�e|�
#��Y�.�<�Ze���ʹ�����hQ��З��_mٻ�>��y񆪛�������EF�Fb�W�k�L�[��)���VZ5�%5x��$��h���qeߥ��DY/��jI�2&׊���*3P/y��b�������}�RṰ���uO�t`�,(9�����ր�n�3v��K�Ӑ�A����6����Qg��������i�����>��ߣ�b?Or|"�R�7xެB�:��" $��U1���Lr
�����l�E0بi�ȖG�\�ߔ��7k��+h���x���OMle�/>u(T�]���7���L�+r�;��ƹWj��dZ%iL�����j��W�H���2�H�j����dT=�DrSiN�嶛���b���\+�[}B��l��0�qA�*P:h`^
��*5#���� ��2鮶��x�4~� Q���Jߣ0�a{D"��.t2�ؾZ4�U�O�{H�I��t� �>��bxk�?>#%�NK�����Ų���Kޜ_2p�S�����b}ס�?z&��8�BM"K�N��xݑQ��m�ֆ�a��8S�������f��v:VW͙���:.�f�T�{^�>��5�H�|�i����
�;��o
s˅�� �ѓ(&��yL��.;��|�2Н�LP��>��kl#b#[sc����\a�m�ꇽ�.�x[��W��hӝ�s#��?peO��m�k�l�L$�P�ٳ"6���6��x�J��j����I*N`�[-�V�7ܷJ��W$�f�'���\ 7��
E�0�^'��Nq�;R��r��Q�u���d�k���}C(�l\�l��o�i��4��9���k�Z��� ��Lvh�l�K����Ou��d�����Iz��4D��9�3�ș�E�AiZ_�RGnAB��L)�7�y35������7�Xx��H6nGP�*0d�_��e��`�����>��ᔌ'�`��p��v2���E�D�4}6�#nR@�R�:xW�+��D�����	_f*5������C����Q)ٳ�.�� ��7�4K`�ل��y^>8T����ѹ5�����)f:�������D:E����8f2�d�z������k�}}v��kH�.���o�V�#~�����&/
:,~_?��Y�����q^`�-W�) �R'5�SFѲ���Dy
${�A�����}e	2�rm�Uզ(x�[I�X)A�4��JՑ6�#6�W�z�RK��L�W����ޥ*_��G�y�3�����h>������:GZ~�z��n^��\0���K��L�8��m̪@�3��
���1��
�`���<�& �/1�e��y���L7����X���)�A��WP�Q��Z�*���&��(=��lq����p[#�O^:eٶ�[��ʡ=ʁq�Q8
p噎)��`�3�v@v=�k��� X?��vI�q��8����7�U�:$S"Nk
�Ri�9}���[�B����Y�cΥ�u왺�>�Z#G�ԅ�-�7�\�h�'7r��U������ �����_��`$�!c\��n��?�'�'�A�+��j�|;�P]Z�a%��#��a���>�K\�9(�:��٢� ��L�[_�U�ԭ�u��c�C�WPxR���h'�ߊRQ#s��B��/�dHe6.�Ո!ُj�΋-�~�NL
o^�m"��
ߪ���W8Q���,6���ur���q΍!qtR�PFA��x���a�ӎ�8�\G'f iP
6�����q�Ng-�{�dn���<rt�l�C����BP3Z����b���:�B�N��sQ�Ksw��g��� d�(?܈�5�2�Ő��b�,�_������в�9�<��ղK����{�J7�ɲ��E)?���s%�o�*���!朋&��|̑V�fdVv�#�R�n�Ⱥ�k�m�e�1g���ʽ:EJ�:T/7�څ��>�u_b�SU%�Q��'x�\��ĕ�)�<c��4�㗐���3�Aϰ�@ �CXy��k�ŕÂBd�����|I�)��]a؂�;ϖ�6=8�������ʞ�l�4nJ�wSVh��	���������z��o1*I��}�DH-�sp�R��m)xJ a�����ap���+Ɖ�qG<4��A�Z\pIKB�e�<\`���N���h�i�l�~�V��6J���N��C����[4H�ˈE��Z}¸���4P�,p�Mrr"O�O�N��v��93��A�x�^3�5D�~9?����*L=��|�l'�wF�o���$U����4L�0X'F̳DnȠ"wt7��.L4����$��ۦ��k�eW��{+5�HB?��jc���$k2E�����XH�o�a|�=\ڹ��X&dx�q��<B��i?��	%�j�ئ�VP-(�����2� '+g�u���e$�w�Wo,{�Yz�U|J�B�8���}�����Fg�����C6�)SD�O�(��_��3�"��8 >�y��]E�&ݍsn��s�L4!�͸���Sc �=�@`����6Fl~m�r��AY����\)��|��}dq�6	�`O��m�`�����v�O���D��4]\�O%�h��[��a�c��,����w�S��!�'cJ�۩j�ѓ:��Q`*�� 6)$>f����X#����� f�Ҡ���;���;��7�m�+�،K��l�������S��Lש�j����ݳ��>����&�ife͆���F=�#��5u��mX~���
�U\\n�ީЖ"O/�+0
�>��4�X �%�p��}FΠ����f>�d)s~�B��#�a-E������y�&s���tj����к���9B���9۝m�(�w�����̡:B��ᖖ���6}t�� �2�R��22 �Q��Ƨ�zG�[�̗�@�?��z`�W�?��&�l�"lYsY�$ϴ1���[D�C?�1�>�����_��p#�A�cn*z�`r�x�����F�;_M�oe<����O�=�F�_�F�M�8p�As��s�EP���2��j�UT$}踙EN�i��]m�aW� [O��`���)d/�{��S�
Y�� X��M
�<�k7�P���|��i�����1���"�m�_��%-���CMy�;��"0�/P������%TrP�/�s3�/�kl%�-�� ����=;*P�9I��f/������#�	;��l3Ҥ#+֢ڐ_�F����TK�tY�L��zo�c�x6�e�Zg6�TT�}�i��������H�o� B&E�(�Q�~�����桿6�W(ZI�%x�����q�l9 �����
=���� �T�24���i��'�A#��)T}]�� 8�1��/�[�\�>�w�@�%����::�n�V�9������U�T�c՛�ϐ����' ��:�]40Q��,=��o?UI�v�?�4,x1n� ���=*��	fP���Fj|PCo�4 �r�IV͙k����������Q־jh6��{�AM�����R��(��G��.e��s�L��P��h8��	���&���SEņu
id�V����w�/<e��8�'�qf%ם	��W��s�2�\2���v1]�S
��[��q�:��za�x~�[��Υ��	]��6"(g�ݬ7~��Q�D�u7e����\O_i�,G�e�a��_�Y�~9�M����n'x�#��Ȥ[X-&��x}�I��*s��m^�ܴ�q�@��n�D	�PU~I@dM�E����I����M�T�W�m�p�����!U=���~��s~��(	�.gn��m������J�-b�7�H��u�v�Yx�/����B�<����3�yvmf��2dqMt�d,	�C�.� |�5mZf�@�B�����p�+#D���;� w�Ew��:����qe��T@g8����b���􆶇�O���v0b9A��!R��=s�J�^�7���&`���!Y,�iQj1!�=]�Ҫ��