��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� rā�SZ )����C.��&0C]�-��[�3�-���+��պݣ�k�J�vo`�A�����f����u�X���v�=�а���]Q�Wۿ�߸�=_Q�X����j>��Zw�K��SvX��ƥ.���#�����Z�0���#7{��\S$��@1I�QX~TQ�E��db����۰� ���>0�%�9�j汈��}��1� ��2���h�G��SeY�a���	'<x�p��k�H`�H�j^y�0�s�78+���ֳ�`�R3dW��_��{p[�?$�s0��#�zS�_��bH
�c�p�IL7]� |����Q�� ��Rr���=��E즕2%�����`�^��l�q-�]�p��jf��Ӽ-f%H���ȳ�>��+���M�71��4_�) 3�46h�rb�J�W� k�h~K0�>P$�_n)���5�r�j��W�J&޴o��$>��6��ŀ�;A~<6P��K�~��f��*I
�Z��}`q���ApC��n���g���3��-�іrO�mF���,�$��@�BI�q�}��Ȥ֐����î�䂧��@������U���vU������ �T#K@f�㯁����|95<@���+�-�)�����K���FI�k���*@�m&���
���ma1[�2�u�I�\�U�yu���o�|��2����;�W�W�}P�K>%5�'�8���׫=����k��,�t�M�0�8]q3���N���GvZ�i�+ C�e
��Ќ�S�v<%���q��e_��
�k�夞��>ZO7E~��5k�TW Aod��eE���G���ɑ-'���?�G$����ќ����8ɸ+ 5ʗ���l�d��,�J�
�^�3b,�����J����#n�zK����z�&��;|�\�^���'e�W�����">�w*	FO��3��ȗ��x9�����a��r����|��)�h ��2Fb��)\ZIV�"/��=8��
ǭ�eKKU4.AE��j����C_G�H7�m��q�SH'�J��� �j�[�'�R�����y�Ιm]�"�#�'��*�~�������K)�r4q�ݝ�R)3���YlP���L����R���m���:��1� ]��p�1����(�<.�������;��=V�
��>[o��}��=XQJU��
(�{4O�qri�a������$kG(=�	O��wu���|��-�l�9Zߓa3P�֕�h���kf�h�� @�Z�z{��ϯ����[:�¥ �Lɹ<`4�W�L�U����,Q@��"*b�i��D�)�ɢ�Ӭ��{����}{[� ���ٶ/ "�T�f��_�|w*�����l�60P�=��5hN1��F^񹄥����&�%��:�����ֻ���y�4�͍��ɿ>�!M�$>��8,-a��O�p�~ �9:�0j��n����V˦X�I�b!�MƝ�^�Ǎ�֗,ƹ8䈭�v�0�Q�&g��1	V�E]O�/��k�eRQ�1����TT�?x��Y�l�g}�2#��1�/��u��E��u��[�<Im�=M��,���MÎ��*�����ϡ0��>���~���^�Lҵ+��q*��x�xf��p�fc�)
 �8�B��Ru��XƘ�-0�F$�E�	A6#@�/��f�pe35.�4�(Z�T�����oG��������>&���5^M�5�!f��X�����Kj�����F�#%,i���3��C�/����3ml!m�:��*J�]�������x4�&�*��Qz~��X ����#�?�˹��J�Vq+�-�D�t��`:P:��lr�SS�5�5	u�U�U_����+�V1M�?@�(AN;�}�O���
[s��h�y�(�����I�f����$�����o/det`�6��է��C �1d��=�k0^*����A��}�U.�d�'_���D���Q`��˵���uQm����t|�:v�������h�}��`Å�`4㒽�8l�97$���
y��9##��3�}ż�<�s$�Ur�_s���8�0�4pV��h[&�,�Ȧ��ð�v�i�q��eBx�
i�	P����x�C0W>A{�d��H��/8��.Xr�jC����f��n��^Sɹ��@~)�<5v��=uE=	��ҙzM+d��¥��J�&=t�W�\�;V7�%��\Q�J���2��o�l)���}�b�M�7���}�}\g�-�ٿ��m�&�Ҿc��~�Kt�?p�f3���Z�������3����Rrc���c��M	��f��'^2�	E��4�a�$X�m�h�U��/��.�l�M��oA�q曢��`�O^]���T� pt�qߚ��o}b3����*Z����R�j~��Ͷ�ʠ/p_C�~[D���r���k0`�MzI*+�K �i˯a��Ĥ|���al�ր�"����?vo��$��+dp����� `�@*n��<xVudE��y�Y�ے�j�gגkN�ʏ��g�	������?��>��N�z��Y�����h��E��muT�¨I�ii�V�m�p1@)�+�h�dS����('��)u&�7Wdڷ&��k��b�F��̱���`�jmΑ��T��M�X����᪝��R(��ޅ��������'�2;����R�=�����K���q�~���|��� �EQ�%��wi��HY,�%�.��e#!��"����+�Y��i���^R`[W'ԇn�N�G֓'��c��([���d�_1�uѺփO{�%I�;��a�
7�m��A��bU������E��~���܌�F�
���Ǉ�ϥ�;F�F��6_g��Vꃩ���/����̽��3���w�ۗ��'�>��N�d�߅)��]�� �C-����ۢN�{e�a�LVm�����wP��yNT0Ee�@��i!��������e���@��걱�̓ݲ�
�86_:����;�!�t�� �n�5�W6�V$�g3���`V�=��:��os�;�H}�-s�ǜڋ�p��m��O�#��=S0�]GZ�?���f~��������5�t�ٍ)(������T?m�ƾ�s��u�%����a�2�'M�)%)�P���lx� ���2Hm%AՄpض