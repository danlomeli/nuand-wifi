��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$��7�4��L+Q���+2�"H�������v�ao4��	�u��=��d=�>�iV�f��l0�Zs��7���~rM��U�`���e����K%�u��ݒ-� rā�SZ )����C.��&0C]�-��[�3�-���+��պݣ�k�J�vo`�A�����f����u�X���v�=�а���]Q�Wۿ�߸�=_Q�X����j>��Zw�K��SvX��ƥ.���#�����Z�0���#7{��\S$��@1I�QX~TQ�E��db����۰� ���>0�%�9�j汈��}��1� ��2���h�G��SeY�a���	'<x�p��k�H`�H�j^y�0�s�78+���ֳ�`�R3dW��_��{p[�?$�s0��#�zS�_��bH
�c�p�IL7]� |����Q�� ��Rr���=��E즕2%�����`�^��l�q-�]�p��jf��Ӽ-f%H���ȳ�>��+���M�71��4_�) 3�46h�rb�J�W� k�h~K0�>P$�_n)���5�r�j��W�J&޴o��$>��6��ŀ�;A~<6P��K�~��f��*I
�Z��}`q���ApC��n���g���3��-�іrO�mF���,�$��@�BI�q�}��Ȥ֐����î�䂧��@������U���vU������ �T#K@f�㯁����|95<@���+�-�)�����K���FI�k���*@�m&���
���ma1[�2�u�I�\�U�yu���o�|��2����;�W�W�}P�K>%5�'�8���׫=����k��,�t�M�0�8]q3���N���GvZ�i�+ C�e
��Ќ�S�v<%���q��e_��
�k�夞��>ZO7E~��5k�TW Aod��eE���G���ɑ-'���?�G$����ќ����8ɸ+ 5ʗ���l�d��,�J�
�^�3b,�����J����#n�zK����z�&��;|�\�^���'e�W�����">�w*<���=�O�V������0g�R��6:[R5
?�b���Đ������ʊd������Y�Pȍb��w�p'~J����썻UZk��+9H3~m}�磌�LOH��b�q)Hy��~��*���L��=G�UZ5�	�Ҡ&8f�|�p@ɋV�KD=�;{���p���d���<�-q0�;�J坧��U�� Ӳ�E|ٮ*���UǏ[SND��I[Q�Z��|�o�Ht0����������/�7�[�R��y��6��5��4��pvV��C'$�����_T�p�Pe��.��D?Y�_��>�#q�F9Uۣ��:�c哤�H�2K�#B�g5���]a�2�~�z����guh��vϻ�N����\1��+jS�%�Uqc9g�,qH�����'q���h���F�)��/fG���XX���žDV��|�6�Jb^9b.�o��ϗ�ek�aIh#+��	_�r%&�z#u��d��~�ϵ���Qwݙ���ԪB�r�X�.s�����̋|=���YI�lI,�f�GS��i�P\�M7���0����v��"
T6�C�+K� ����Q����Rvq��ʬ$��\�+,���kߛ��!�k���$�L�(���0r/�I��������u��F��$��=jFG25��w,����
sU�j�6�{=�T`�2؛�@(T�m�U��5,�����y���S�h���N��*��#�|Q��U�&]�T�Q�4CI�iY��g�'�l�6O�B�K�{`Sۖ�@�����V�W'�A.��:��J�O˰��([|4�o�����	_�Y��ōS����^���Fy��_A�M�m��_ϙ�`"��N@���,�r�D���4k�������꜀�ퟀC������"�##1�v�s� Y����F�ޛ/o:�'x뻖�)@F��ڽUA����Hĺ������u��h�1���k����FɈl57c�]t�Vѵ7�N�K����,�q}5�*i�3��J<Vsk*Ő�ךc�M@0mw�GK���'�ȚBe�#�"�x�7�@BMݨr:�[��� ��
R��7Ъ܄��v��#���J��5�4��Hޘ��P��H{��o��F{�4�{�{r��#���Hţ,wG�;�0�*�9�CWZi�s�J� e�u��j�L����_�D�9s�)�}��{F��馿7���`/:ÈD�ZWμ/i|2����aHRGX=�(���64kC��lDrI�:3���,�!�K�P��9W�*��n@O؁��)����S������}y���Z��z��n�L����G,����2��R�	��n6���%Q�!x��zi�x�Q�R�S8�f� �A[l��*����#������_}���{�lsF���]��ʉEV�!VO/6G�����6�Ǉ(����H��SMl��a���f[���c��F7+��6�m����JW2�@J��$MߐhY�w(%��Q�kܪ>��7���|*oVx�Ȍ���[+�"k�Fb�e1��XSm�����.��O|��������H�1':�� ֏�N��֤j[_� {����W-�����m��*�Hd��B���O��;}a�0� wgu�1����J���d*ȲeH��A[�.dbĆ,�
�Ŧ<G(����\ɧ��P�%/��.���2�e��]X:v
��^'���Z�a����T�TG?���r�e�Qt��ƀ��5
�jZ{˨k�m"ѳ��_x����'��-o ��my����g?kHLOݥ�!E޺ȭ�����K�~s�a$�5�}]T�-r��N,��O�c�c*��Y�\-?7a��n���p��2��*[Y�N}���f��L�m��z=��"�(�/�����f97��io��L�8�AY�Z_�.:=�g���q����ٿ��O
4�O̅K:�
�>�w	x���q�O�Q�-�)�yb��;K�Һ�ڋ��Y'�R�m���jRj�Q�
�{������,�z**i�_p�=�+oG�=%a��Ն�V�X8`�\d�����+9��IE@2-���ñ%6!�〶�?�0#�kGPs<]"f�B��tt�����g_�R�&3���=y[A+����ix-�%<�N�4W[��������s�n�����H��33�o��_E���z�KLl���l/U�M��=��O�!+ �d��v�R�D��W��C<s$7V������H+�Fd���
�(X�M�"TK����Y���$� ��;��,F���+V� h@�*Ѕ��T�`�ݺ�B_�jYt�����ȘD9D�o�d���t����u�*=x{��	#����:y`h��O���n�!�dN9($�~�'ý�{�B;Cu��U��V�*ʷ��c��g��f��)[��dSy!���7pw����Zy�عl�I��mZ����o��]98X�[]���v��g���[ʕlpQLi@�u3�Z9[�=y�=}�/�WUf]��o7��	5�V��ۈ�J1I�ڕ1k�[]��P�K���\�dlFI�c�.��tcD� 9��T���=V�BK��G�5&r�#�u��|��ǹ|=��w2�|E?�T[��.��~]��NrC�s��q������Zd��9�LS����#�O'~cǚ���5��#籝:�I�C�˅��xu��mX�����Z�3j(3|�M��3�N�˴�kFM���,��)*�N�5T��C�x�Ԁ�lq�((9�t�TVr��c5`����к���'k�҃A6�~\&E�q?���|�(�T�mTߢ������[���d��˖�t��|>n�=L��=<�B�q*������)"�	O�ӰW��#�}Y,�b�M9d�����X��О�3�c~^{p��-3��ismz��2Jq�l��z�l#�e�& "�*;����~$u}���I��k���C����	%Чï����9�,\�L5oA�f��*�p^�*x­՘YD\5.��S�ϫ' h���|oVxtTk���i>Ӝ(|�2���F�F���yD��j}���em�����s��t�({��f�Xg̥C�Gg��'�G�������yF��͞:��Kk���J�����$�d�ɘ�?��.��/���"i��C>��YD�[&�F*�aU�nN�(oZZc�%߅��HIMB����G�����Ε�H%3��QC4v;�-�B"�ﵦA�����oR��W�dZ�8G�f1������)x���"��p9�*Zl�ᎈ�%�A��?�mq©�yH�����Y��Ke��!
�D�@
��5��x�����n�[�a�C^����iLEb|K&6j��u�kX��b��x���C�W8I��ղ�t�L����B�����%�!����:a���^�"�ւ�]�L��匆JyB���\ �[�_�4��_��z	t��*O�S�כaA�t^��$��픰��c�'f��A^���O�q �ƩA�� u��|�;�L.�Gf@�ץ��w���9�,�3i��r=�T�
��0ʉ�ge
7��wbI�7�Uwb��:��>4��Nlɬ^�c���=�n8���M� �Ժ,n�U�&��#�d�� jt���Ǌe�.�|����}"���n�0�����h���d�D�#�R���5�>R;�������9��z���Pb�R��<|��^�7�e��B�������C12�F�{�AJ���tf^Ya�a� �V'���,�J�'���3�$ �t�9�+#��|튩�l�'"�]�����-���t;ߺ�<Q�AJ<��Y�#�+�ٽ�|����H�;ׄ�[\�o,Q"MKW�3�V��=&��7U�B7a���|D\^\�`ʁƥ�b� vy�A�z-4(��.���@�?<�w�C�Ǎo!Kos5v��w?ԃFȹ�������ե��|3�\���y�u�D�8����ST��
ZF������u�%��:��_��BW'Fy�	�6ծ��7od�3۸��{Z�;�+L���v�"���_t.�"uĖ���a���þ��R�V�WG�o�\����@sJ�իjY�Vz���=�bkؚJ��WsJ�o�&� �5!$���[��M9N_�����H�5O(Ϳ`����K��$�1G�E��`�`0���'�� V��do�D�)p�� �'��l�V���g윁>5���L.�E��X�5N���M��6aYu�K�c^�`]N��i��:����S�Պt��"~2#-̦��Z�^n�dV�0��Ͼ>�oj��Sn�0�Un6L�'aQ�Eoj��<��6��:'l��k�+hU
��� �v�0��U@TI��r�F�4����i����8(|z�s�r~�<�J��3J�7��n��&�T���'o�X����Es�K1T�
e1�9�*y	����ހIh{c�L��)P�FV"�A1��1=��<��qkB- 0-!tG��6�rjn.T9���n����u�� P�D��#��>�*�^Yf�5��kV7���G��-��������n����Q��q�0�~��z9Y �T�F5V�Uʡ���+����0��^��&7���D�LK�kY��� �T�Y�IA��&&S���l���d��Ui���\+���f�#���"N�e�owb���V��	^`6��ᚣ6I�郰neF��NeԸ��H��w��e��qQz�>��=H���(��{�9u-c���h��y��8��Z�V$L��^R��qU���o�����#� ��3cR�4𺖮�A:�$7����}��P�z�4��a�퇡��ˣ�a��]�_>�����^\U��wX��p!$(�}9X2��3�ǆ>�Z�'�
����O걹�H�����<��)9Q���d����� ُso�	�M��`�Sb.�b�~θ�CLǍ=���7y^�ݠ䂧�*^�b�?�'� b����Af��~b��>���z�|w��f��gI�9P�Ŏ�.'y��gs���#ELO�c�b�w��y3��hݘ*�)]sM��1n�� �B��;-�<�:�:�:�/�Tpv"�:�o�Vh@!�4t�P�Gy1{��S֞ �R�>��G�8t9V���	`q[%�31�j�9J��;�����V4�}�`x"�(��(��
4ElR%ISqa$"�?O
�<ŉ-E�B%G��{O�"42�
�ÞS���
V<����/�uhz���4}�N�`�@��l/ŕ� �RUcS���PQSܑ�D�'K�S�'��R��^�� Y�w)L��MN�a���ʰ=��o�
9�#6 xi6��
���/��Þ)�5xS8��)�<�\q(������w��J��+�L�g[��⥀A��;'7MFi�g��fl �v)[F�S��/�Y�Nq�jڄ�Tv�yZ��o��:�m�ە�n��)}�=����l� fڷ9?ȚǄ����G,��Wwf���7>N���R?�V�����F?���{<�*d��(¨��V�$H!R���6�\	4�u8T�}�>���@���Q	�;v(TT/�y���ִ`���z[t�� gDߤ��Vm�͙j��Z4D�����P(�O��u�
p�����f�Z�)>ܖ�sPBh⍿8q(�Wm���[o���UU���=�Z@���R8�:�! R.<�]~���<&$�S��h�E#fN\t�����mP^�ܔG�?�)�N�C3�p����rw�x�F�t-���:A/OH��X�۷�fe����LM\1-4N�����B�7b���Sy���L]���%mwR��׵@��&��??����.�/z�I�Ξƴ�q80�Yv��L8�3�QQ��l�E_F� P"�U�rF�jt��G`����d9����i�>z��7�p�V�U!�`<��0[>ڕ�G�F������v���>Ƴ���P�ݵ�����α��$8w:�O�?VD�0C��b*L� �Rm�P�PTB�f7m�繄~n�z�׶�n�!�1��+Ewz�᫥�*gB���Or��C(�ד�#;����kl3�o���Ծ������.�Gߞ7�&~&#�H<��G�-n��$��u����8;�?Ak1}ly�E�;'��+�c��q��W�:�6��U#	�ٴH������K�$�ł��C�\`E�6�I�.�6K+vE�.��q$�U�A��3�Tr�����_*�������G�'mZP��]�@d�%��RR:�	���rӮ1���n��w��KZ��N0�>��'Q0"
����Ɋ���
jL�?���K��_K�tJ�__�/ڶ�C�|.+��\[g�}Z��4ʧ
@���|��A�����G�m��~���. 3s���_E����v�)�>����
�$�V��w9��ĕ�?<����K6ݝ�1����^�;;r�x��8���!�������^]	��7,�_Eӧy����@n��dp	�/�ͼ�y"'�=`����d�VFC.m�b�-"�4��o-6*6����_`�!�0S��Z�w������O�`�1o1�ū��X#���CY�י�zɨʟx�e��g�bK�tǤ�	��O�ֿ�mH�0Ϲ2t0�����j�;5�yO�ﰃ��<��M�lx��j�
\:Y�OŸ�'ڛ�)2T�+v�[�5���9rU��T�x��ӀT����1$�yAFy?_�2\]�XS�*�w:-k�C,
�6G�hp�Q�.�T�$��R��)��onș�z͸r��k�H@�����bZ��� #5��8=#cG��L�K�j������o�ܤ$T�IP<��e��>�Y��c
�h�ЂݠI�+A�_T�&gq��-K!A��k�����A�Ŕ��|&���f>�,n���t������#�Ua`&ޜI�(���ʨ�j&��+�I�6U�pu�!����	�hX�#-x�21�ғE4��ͼǅ�Ӗ���;=�ٍͻ�����Ɵ��
eqIc�A��G�0�ӡ�?�*ߤ�/�v�G.	ֵ�	��b$�b|6������=5ϩ(5�2�f6�ZlZ��A]�ZB�mG���I8���?��O�+2�/��0�Eb�،X�2��q����^�����F$�b��+����#�H����ir��#��uU�2�}t���W�1#�me���1.���0�%����gz�y{ӳ�Vi����l[T��+���������zd�߈"Vo�v��eB�[s�fܑ�%'��'��Z*'�#�_�4���[x��k�o�e��g�ڥH���g*�����  �[�^H�i��:��������Y^t	�Hh��#6��j�As��W�i̇ef���dź�5�l��n�"�K9O�F�笱�}ѕ�����=�Ȁ�?��4Χ`��4�Z�[p����u�<D,�2ޯ�7��5re$��3'�n ��Hr��ʟ!5��~jy�<�t��ٷ�y�kȾ���H%Z �),iZCb��u��p�{$#E��W�ra�;�����v�<���Q��x�����lN�¢&g�{��Zv�uNhi�G�~�a���}�n/�Ó&��<,�����x����୿�K���V����
 D*UV��L]?$`��J��@[��K��l	2c�i�nZ���M�>U�N~��)��4{ϛ��J�[*;��`���J�@�I]s�奧0�U���Q{�/�T�?#���W%�G�@�����%9�.�GCb��d��	�8ƙ@��l?/5J~�%(܋��A47L�
�^�Yk�{R%�NQ�<�[I"��)�*�t��a��'�~�YO�Do"���<��i�l��j���\��H6�Ƴ'4��Aդ�҇��8���]}e�`�\��Fޏ��}�QC�4����J���NL-9��}���k���F��_�4��17�e��
����h�V�9>I5�2[F_#9g����Y&E�C4T����x�|�	Bp�Ք��e����7=��^��YX/[ro5��/�{\�!���T,$o#�\�Xd� �w����~x:iNL�u7�Т3�XP�j-�j��/�Q����(/Y (�.�����V���$P\�
�k�@e�h|9c�g4�P��_�+!d�,�5^���G���tbl�<�����a�O$�(X;%��HI>3�dq��m��Q╔��l�M�!ه�e�_���{�,��=�/+�}cJ�A�D�;�+�}B\I�F���`�e�W@]@�������B��t��\L���B�G�n�
�P̻���Ӳ/�l�;Q���x]�fM;u?n�Ȣ�� �xy���]������ �a�6�i� g��a��Z�m�j"u,/Jʷ�9�|Z�	c�I��Ԓ�����76��&�$nS���@,!��d ��c��k{�����@�cć ��&��M�v�h�j�N9�b+q�D��T#��<�b�Iq��6��w��Ls�\��9���j�/�q4�-܂c|�Y�ZY]ts/��3v���Q��P�~�'�~�� ;I����3o�?�4�Y٬az��:�0��h��G��\��K^;HBe#�D�`���h�	`�R]����a�y
�O�S�	�oۍ�z��cH��V��9�D�#=xr�R)���>dlh3D6m�b�7���e�6N�h���;�@�S���!ό��r�eg�d���eX��ݛ^&��UD޻L(A�� ��׭W �s*J@�|�'��ڶ8���A���bl�����_E��m�O��8z7KK2�@�>���ù���/C71U���V{|�f���X@����`�P[��jL@�,+cu�&�/C���l���vmE�bp$���w�D�#�o��D�H�����W��&q)�e{^�%}��\ꏠ�;�Ȋ�׸���gBy��׬���I<�5$\��td�K���D�Ƈq�{ot��f���V��g��>���ix��0���0Ǘ(��@B�����h��u�G����a��`�^�C��$��>�6ԁ_Dc��E��0�wC��:|5@��cO�L@ڒ7SP�`ݽ�!�m�bp`�X����S�����7(���:��ne$�/��W�;��Ӛ{�(�$���s��o�!0��i��Qa|ޱwIH��^Ou݇� I�5��邀�>_9������{�rg�<	�|k g�W_b����[FN��z:�Y��QI��MLȃ��ɩ����\��'VK.��V(w"��s��iE��(Ą���t&��%݄#Yj���,�.���ٳo0��.ùu/
�3z��x	`�
��M�sil�Y�G�	�%P�F%��ի4̚��#H��8V� Jw嶌��gE��,�n��Fx�$�I�)oKqi����S�� Aɹ�0_o�ZF�ݙ|���)����2��"U�G�H�O� ���7���r�=&@6�5�@�
�[֤t�����R�_�L�g^��-�E��3�/bܔ���^I�� ���j�o)�QMn$oV��;zh��́1֮D���=���5��5d����|�x��#�u��I<�CG;���P��:��7�<B��\6"/����җ�����������c����\�P�0�Χ��xxY_���e��85�K�ѱ����!b.Әqu�"֌8u��RL�GOg�Z�!k�� �6����I�S��CpUn� ������S���n���֘36�$� ,r��4ks�D����F	�����H�rb����j 4_��M���,~�b�	:j���QkFBsұ\)�Y����*4>���)o=B��x�6��޿��T�]�nLGy�.>'��D� _CU�!F����W8֪6S(Ò�h�#|�9�jA�2��4��ʑX���-2����⪹y�O9���z��!��_��ruO�'�%�c���/������Eޘ��F:-�|$��t@y�k1�4+~�$BxE�i�� ������"Yf��'�y{�=u)$X�Y�����"K�_H�5Eh�k	��Zn[�������=��G�;~�b�t�����-W]u����
p�+aUA��zV��x��MՂr���0��5�yT�����k@�7Wj�v��*38�ߚ��-GG�y�[�xE�	���O��0��<���p��p���B<Um�H����I�n��;�{��O��u;��L��	f]쓖�ޫ���l:BT3�	1�W�ʏ U��>��/�*X�§����6=.�=�f�5cp%�4$_�x�~��$$�G�Q��g2e����+3�bI�ý~����Ƣ/����i��5*�9�~��ɡ='�)�L��w��=U��ʦq��i�~ڲ���[�Ÿ���P��=Guv����w�Э���_<{�v�*�kA&��9p�~��B8[i���F��*U���e1YT��xs�u��6#
 ��F�&��^`��c���k�j6y��hpPo˂�Ò�U����l�w��h6�C�'�R��n��6S�M&0bV�c�7s����q���ˈ;-z݅���&8�)�d�e�þP��8��0�:�Zf����׮S�D?��`�?2�qt|��j@v�E���5��-+'BJ`��Mɠ��r00�$;,��<w�M8Dd92p ��y��
��w��SU��vR�z�9?�ǽ����f��!�לn4�K����@U_G��?����''1%b)Z���+�^�%崣��O��)���"�N��i*�jC|�8P�х��D\��<w���os|��K��~ �&k��
ϱV�'���9N\$#g�[��h ��H'�Z��N��Hn��#�������[�h�	k�z���s�ִn��&٢.�5o��ӿ��/���s����"l���<�� �{���1>!�u���oY�S��%�F���BZכ[��"C��"�I-����{�����rf_Z�>��[#Pv�?�&L3��}�*��ن��w\��K��`�X8���M���T�:	o�PD�J�L�fʇȀA�$���s4���'�K�NL���r�"^rdb��q���������:�mZ˽G�!�>{���Jޛ�P��1ޑbW;��L�J���zC�K}&2rJ����_��Y[O_�e�;����|D��(�ٕq�i0�&��y|��} c��玈#�Y��3L=�ϭh��[=�؋u�l�%��K�ӔD��$���ϵ5���[�Qf��`(.៍Xr���% Ol�˪-�$�o�I8{�ɐ����m�����Ù=���7�i�<�1[��w����{.�>�!ȡbM ¬NR��z���[@�78����0�ٓ�
����Z�V����j�4��!|�Z�IWc�d���g�;Bc%S�{�"�:A>��9=a�7h��;B���jV�C_��k���]�H!��v��;�ܝ�a�;������>�n�.��i�:u;����+pV��U���5�{u����$+�Y��4d-��M��)CJ�<XS���C�@>�	Y�1H L�)�zL}�t�)���&��a��� � ����>��5�����O��`�zr(H��'�+��qD�O�}>D��/F���Ï� akM�Xc��!h��lj�tNdP�nav����|8��(;���M>3c�)���#%}b�)�v ���ج�݊(�u{�^,9빳�����3�8	��]��/F�gc ����"��s^u��\��H���9�_�� ��;�5\?��T��L6�6�P"�%I�����H���ָ�T] 0��[h�w��a�u�-��)�~q����t���@�4�����d�J����l��Q�_nT�Y��#�tj�$������ �I��:Ѡ�bۄ���a��N�;`~��杗nA%�r
�?�A��z��{� �Q�G�P�"@CF��[��ڴ�ꋇ_ߐQ�"��݂�tYm�r�������ŕE�PҬ�uȗ���)�z��@<46QE? �·�����kj����r�P�
~]/	s������	>z�ֲ1��������O%!<D����*@+�A�'w�NKn& ��1&|#���Z\���z��b�ojb{��j�I��`�r7��#4{�]o�L,�#��~���R�~;��χ���x��vR^�,^�~t�۾�6��/��e��Ӫ8�����%�y ��	�$��I\#)��xbfU#P�[�cW0����q�\⅒��{��|**����R�Ӟ�+p�c��}nɅ��M���H=H����������b��{T��
�3�xݾ�h4�+�:�~~�[N�`���<D&� W/��g��<U�<�N2̗ ���Ʀ4T���h�1ǣ4_;3ń��}�Á��\��4s�tx)�>8_�=�\/��+�@.�mB+�k$�d��1~�=6:���QDd�2����%�]���?�`�����V͈�s�P���Zc�y���].�ޝ����
~>��X���4�Ia1�c�H�4����EF��D�۝@R0��;��j`"6qM����EM�9&.{4+J�fVm���saG���!nB:�������pGA��Vs���4�د̇��,ׇK��p	��9�˟�;+�+l����	\dnI����T�{�@ik�� �n K\lc	%Q2�3:�J������@��_�O�B{�	��Q������H��	��8F���`�Ӳ�=�9��b_e��$�d����`t1&²Ր[��o���a
)PS���ʥ�tWAh�B6"����;0�ĉ���}�q��U(l���B
"*�bbNfZ�}yNc:\��1���f����ν�������D�|�.Zg��p@A�w	���56����#�1�I~�4\2�gtHd�!�-���Y���0jt���wA�F�ڎ �X��5.e�MM1�w�B��l+��v����>��9��ߢ;��� �N�E��O-~�^������*,�$(��S�}�Oh�耍�n�E�x��Љ��w�z1�C,�/Y����z�IA����T�2/�Ǝz�y$����c.��,Y��@@'�&�|>�,�J%��b�����8�̿�������!��DH Șm��UA�h^�x,v���T��U!�b��E?�M��qQT�����pZ��	,	��V���-J��M�(7W�y3��;î�Q���x}���c�o{�z�,�+t�)�����:E��jA� ��8�*�G����E�'t���Nb�>yh�m�;��yʱ��h�a�1F�Y�넼#iJ?��d��lꄄ˟/Ux����8)?�� Ak/`�ٗ���tf�h7�g��m	v�@���F�J���q��	�h����as�CY:Y������V��W7�@Ƣ�1���om��_ݥ�TРY�X�df�K8�ON�3��պ���W5��0�`��R�(hGѠ&Ȕn*��J[��D�z���!>�6#"�"��>2@�E�%F��о 7�s��Q�������W���f6�	���A̬���s�������l��SC����˳�x1"z8T'����)��M�N�ͱ�7X�A�r��> ����YJ�:`�s!��4��x)]�:�6ӄ��_����@A'9��
3T�r,�td�5�ܪdp��t4�z�0��X�cL�I�/s�\�?J�y�p��D��bY	���D�Z�"@��CJL\�Q\7�r�G�¼C�+q�ߕԡI�`WD5�Y�ZoV{�({'ϥ���=_��
Qʍ���F��M�0K��$���M��wrʓG�ՙ�`�0#=��N'x&\��s �B������*}<=���m�v�䁉ç���8�1��|�ˢ-�	�><�%.k�@8�M��ok<�eLz����G3�<9�FE'n�b<�����R$I���l<c9��FB�{��Q���=�3L4��p�0�8��Yo��F�t�>��:FRv�\D�1҄�*�XDX��rb��:����wo�B�=ߪ��j�C���5:�oA����c��FH@kf�����JB��}��$�2���K+�!VY��;#� ���ݵ�m'��$��m]$���R�:�&�˜DZ�%�%��5�u�=T��d�&�l�C,� �N%!:$�r�B��zA���R6Ӷs���b�����-I�.H����_�r��q寮�h��|@Ʀ�������gJ����ko#2W���9Z���.�@��*��X�7ԇw߄�a��S�S��\�D�t��B�1��y�p�	9�9'ݞ�K
��\{~ّ�Ҥ��6K����T�i�o/H)/]��_i[�\�d��7A�I�o�-~��E�?r���1I,Oe�d���$�=��ǣ�i&Sw�����X~ǉ���l��ë.��vӈ�z#�P��#�bN-_#u��6g����f{��_]�/߈R0�Y6}��Jn]���k��1Ԥa���HXpq�	�f(Q����9����M*�/�|u�7^ktBO?eth�T��6M����c.��<cuԜ7�������:��\�c�ڙN%\H"7���oHvğ&�����t����e��;��S��wIJ�G�!;OPtŇ8=��&--��C��):�{�����(/O҄.�0G��S.W�>7`��ŋX+V�*����(���m�$_��{D6�M9��d��L���I��]f&Mf�{(� �,0��Zٍ7�E(mK,��%л�n#�Вп5�����@Ӕ�A�Mg�'�zݦUA�""8u�W�E��H��:���:�a�4&i��	Ε�}�eg9��Y����]�':����d�
�N
�t�(d�K�,Z��+� �x� ��謢K��)��Z�@?,{^�sm�AEʳvgnF�"!��Z�?�9:/I�fS����A��)o~�I ��Kt����q!�~�%��<��;��P>�́O_��S��(�	̃�ڐ�k����%����f��xIS�)pYh��U���tH�1�v8�f��pu���n9�gam��DSb��-]W{"T��m�������G�o^��߇�� h!�o�%������ǿD�ֿ�~>&��a�j(��Lp��}Zk�kD�!��Ud�#�����þ��V�-N�A�\�IĮ��	,�Y7�$~���i�X�A&.%q�7��ל}t����\<�Ё3�rx��i���+�#�5W�ˁT�b��;&h���@69��`��,�%�ȩ�H��p�01�Vx\8���L���ckx���G�H)U�����[N ��W-XY�i�$�BI��u�sy(i\��*��4�+ٺd��lW����YC�g4mf�,�x�>g���d�62DD��wo���RQ����	=i�vg����8��^E�Z��E����7n�!��`|���DC9��<YU���Q3�3�x@��x�{�6�=��g�<`���T�D�2�)�6j7��Χ��+���O��^Y!J��W$ۃ�TZ-�\~��rxaII^��H�m����ASY�W�u�U��ꔄ�]i���q���GR��nr�n����Ґ�Yȩ� 3���=��p�=���ܾB�2|Ui�#�ߵ+�C�uC���>q͕�z�7S�W<�$]Gٯ-`��4`���yWպ��6+�0]Y� 
�";Ú6���C��ٽ�֎�$x��Kl�9HDu�@_{'E��n��NM�	�sr%���<��{���%%��qixԷùͮ;p?�	�n��e�!�9Zc�x����L�8{��������`Ϭ�~���r�C�Eh��J�3���}��M+ǫ[ю�K���]��Jr� }*8�)�.[�II�j|V߆&$}F�w�����Oz�yu