��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� rā�SZ )����C.��&0C]�-��[�3�-���+��պݣ�k�J�vo`�A�����f����u�X���v�=�а���]Q�Wۿ�߸�=_Q�X����j>��Zw�K��SvX��ƥ.���#�����Z�0���#7{��\S$��@1I�QX~TQ�E��db����۰� ���>0�%�9�j汈��}��1� ��2���h�G��SeY�a���	'<x�p��k�H`�H�j^y�0�s�78+���ֳ�`�R3dW��_��{p[�?$�s0��#�zS�_��bH
�c�p�IL7]� |����Q�� ��Rr���=��E즕2%�����`�^��l�q-�]�p��jf��Ӽ-f%H���ȳ�>��+���M�71��4_�) 3�46h�rb�J�W� k�h~K0�>P$�_n)���5�r�j��W�J&޴o��$>��6��ŀ�;A~<6P��K�~��f��*I
�Z��}`q���ApC��n���g���3��-�іrO�mF���,�$��@�BI�q�}��Ȥ֐����î�䂧��@������U���vU������ �T#K@f�㯁����|95<@���+�-�)�����K���FI�k���*@�m&���
���ma1[�2�u�I�\�U�yu���o�|��2����;�W�W�}P�K>%5�'�8���׫=����k��,�t�M�0�8]q3���N���GvZ�i�+ C�e
��Ќ�S�v<%���q��e_��
�k�夞��>ZO7E~��5k�TW Aod��eE���G���ɑ-'���?�G$����ќ����8ɸ+ 5ʗ���l�d��,�J�
�^�3b,�����J����#n�zK����z�&��;|�\�^���'e�W�����">�w*	FO�Δ��v���I�h����p�=.�vG6(bh�۽��d�Q߽`8"�5�I�I��l��vq��(q�)��b�/2�-A��Ⱥ���%�N�ݙc=�ĺ֟_�V����2d����ʘ�g�����!;)B����:���-��
�����G#�1!���/M�P��<�m�<��ٜ��nE��Æ�4	���V���H3p�5I�C��P�(�����ܔ��,�����gi��f�����8 [5�[���R�@,��S��b$�����i�ѸX��A�F�8����SֿT�S�}��l3�ȭ�)��'����<����\���4�׶T��֍�IN鹏�����}�Z4зe@TP���	~f CAZ�T6."����-�XD�8nG[�c<����zUl9��VC@U��J9�V�Q�LRP��`�U�m�ɘ�#u*Aȶ1����|L�JO�l��I�f(3���S/u�"��N�'(<�ә����ic�ɇ�mjk1�p���Ub����!�Lu����M�����;!���>�75�0q ���6���m[x�,�F�`[ΰNO�I��x�Yf�NM���Q5ȟ��Tp=1������țQ>0�����#����'� a��J�D�� <�令&d�:VuBr+^lᬤi{L��-?x'/lێ�ܞ�����7�JҼ�i��G��7��՚�p)����DT�þ���䚖m���}���=�X�'f�=��i92�y=���/E�z��+�lAd%S�./���j��M7�����W�V��bK�0 �ZR���l�B�WkU%BkӯZ�K9#lG=�j���N{A�7��˓�Mg\�h�a�9�l=4�	~N�Hѭ�m%�d�:�JQʔ/G��dƚ������;�+p��>�ë�7��5FF�(��sY�,�� Η��I��eX���#�W# M\f��;��n�-�G��It�-#b���˺J,{'�����#�����.x2����
�I��\�~�-Yc�;J'&)��ШY�*3�fL�X�{
g{�BSs�e���E/�_l�'�|�,NB��E?�<Q�G���?�X2��G?O��Х4_�JGw�>�G��l�!��
D��h	0`�B%j�'�7�]سf���!��N��c�y�pR�i�4�Ѡ�l�8��V^��@��M�����Z��ɏ������Eyr ���J�E M|uס�n�k��Ec�� VJ���GΥ�i=�=�:򬯋�j{��ɏ�(yg*n��Nh�l�n��y����'�Ѧ�6����Z�{�<��Q�mL���nf��hU��d��oS�}j4����h�\�1�-��d�p��H>=>����~I�B,C����P(���CW��J�=���#k���5�.�7q9Ѩ]���a�Ǌ �.�����R,����w�ص��RV�7��� D��c�a�n�lG\�y''��3�O�,+1z��Z��5R_͋9Xbn���y���߮6c�[��&����P�!�� ��ˍ�lb�gl?��p��aw�X�^C)�E�_�rG ��JJ���i���� ¾Eϴ��c�lB�K�w#V
�D��i�������fXImZ�S3;fQ�=� ��ڬ����M���Ң�5��¯�Q|�"fg�k��{����#o7�2�e�W�g���$�|X�H��!;� D�0��#�F���E`Y�+�s!KF��Spdr<�K<�/"�qfs��{2	�����y���	|�8!�s=%�����z��]���-�@�-ܺq�Y��fS(��L1��%D��&�a2��?34���:���']<񝭥��-]�|
�~Dr�c����f!��W^g(���X"�{md�xے��{߬���u(���ϏL#��释�ˡ��>8[2��ӏ��EQg2J ��Y�.��]$�(��3�߼;,��*�<���?J�%����'�F��E`>�{�6��ӐS�K��?�����!˪��!ކ<���)�s���������R��ޯO���a=��m���v���{_�,k��0����Y*��-3����`1�!�2~�P����40SPѪ�7�3_P�N�K8"o��˂��WI�����ǅ��[�σ7�cU+];��p�5pվ6�D4'F�j�v<�: ��cef�颯oЋ萡R�!9���e�����ʹ���KL�G�{��fz���ߨ�{>�����'=0����"Y��ޞ���`�9�m��iml ����bm�'�ߪ �߅�3ݯ�x|����V_aY�z�y���aT��!$�iQ�!�)���P�Y07kB�/��(yM��"}^���M갛ھ~��̽8��G0�X�(α���+l�udmr8-�A�-�������5s#; {Bl0H�w�e��Ƃ��>�;�RL�bC/''NV�33!D��pU���VU���_$
UTw�)��C��<��qG�W@����Ye��~���n8�Ɋ�1�VV{�=��B����2z�ܾ <R�d{^��^A��2��'�缩�0�Vlr4�|�JA49�a[�l��d0�?�)��Zl���-�!�ȏ.oOG$bJ��~��s#���$�k�%k��r�tׇ�vIn �Sa�7̺���l�֑i��D赁dЄ�����C��<p�f��/�ح9�l1]��ɉ��ik��E��pU��:�a:^�\�nsÁ@�-����޹�}�B yD�N��a>ڝ� ���֧����e�����Cj�5K�5-a�u����t l�=�Bw=lv���?ڭ� �m])��܀�7Q���f���s\i1s�J\px�T�P)�I��� Y��J����^�}��,��b��׺���d�o���	_�-#�O�!�q��G� �l�n�:�FE�EB�n�1P��8yֱ1��;j
w���؍GN킠�z��XeڂۙS�FJP�[�ԣP��Wk��O!���(����of�����s]\2] �\�թm��!RV��"1k�A�v�7�'��-3��_�Zλ����d zb��,h�-�K�p"Ia����P�'����h�_��-��y�p��d���^�a����Uu�c����^���~�ynK�܁�~���=�����D�ZS���'T>n�!s�䕴�L�W���} �Ho=�G��/Z�ݰT���=5_�-[f��5 7Z{�6���T}TȈˤo$��|~�S��C����V�35���#�%��\Dc�j}-����X�L���h���(@�B���2���ݳ<�������I:{߫����a��Ƭ.I�?7�������.p�nTzd�}3$��V��r@v��fA+��d\�]� �ݒP{���1���e�� fÙ+����I�Q]8j����>X%���4�8~�t�P
�i1I.iw�3Ce ��0Vſ�	=��a�6�/��@��'��d'���r`3ȎI�ݓ��A̩�G�+�]O��T
�νS�A�P�揽�Cw�W�8�q��e`:$*ţB��|Fv�ih�� �A��J�u~�\P%S�mw���(ힹ����a�m�� ���Ł|�{�|������8�������<"e�L�rЩ��χ3���Ûz[���G>Bѡ�[]Yc�]����Ov�;2|9�"-M����-�*w�{<4�e��[彭V�����Ҭ�S{��^"cTݧb���\�u�!iw���@2�Vh�(��Y�`����Q�g�
59*�8���r[�X��m�*�PP�{ê��O�v��'uW�rW�϶>H��sUz�$�*1��j��$R��/���DM���B':��,�	n�i0���}���3EY��ܺ��W�Ɗ�������ׄ���j>�6J�;{�^E�	��u4y���b�H�{j	�ć���b�1�ځ>�̮44	-��w���/�վv��Ч	T)O�d7� ��OS�d8>�,�n�����A�2U­c���	�E���z$,��p�zI�A��qf�4�/�!eX���<��l65��sm�М]=��I2�??��d���,�����Y}dg�g�] ǅ�G/���/Ne� �&��a>c �V�6�4���T��xe��L7�tS`�[�v������mn��dw��7הt^3ڏ-�=�M�Dx��G�M�B�l��̚m�E���n
6�Q
��[{d�S�&�T��g�W�:��S��&�mptD�6�V���$0����ݧV�\�����J7������Ʃ'�g�Zﻵ���zz/s���J;���R�A,tAu�wC�Wu�m�'W	�T��>���E���K|������c!q3����7�E��u>�F8Vg�P�U���� ��H? WV g�2U�a�m���p�o��B��xWD;{��lմW�7����pPӟ�%��L0��)�Z���0��veV�p����"��Kǳ1|�8$D>�$�>��Z��'U.ɰ�|���b�R�t3>�;�FAY��JN�q�5���B�~'�ӯD1)J��&T�'N��@@'������>���M:y�͍���C����װڕ���!���u+�zZA��"�6�_����Ce�rt5pe�SiRU�$��\���W\��(�C��O��_���P���@5
"n2�Z��v�Ft���_n�s?�!^{��}���y���������'9i@����K��T�S��+ζ`6�72��T;8����SV�Z%Ϛ����(셊�&w�/%��������?Wa��Yf�;�Mzt��	��"@���;��>�[F��<�U��-d$�-�~NIj�~�@>��K!C?�t��,�+A62��b&OZ?����*oy�qE�ZkV�}���kbg���`to���Z(8���������IAR�J
Z�&�|�YK��	2ض��~P���2� �$��Z<'#�3"���w�!e ��=�<r'7�0�d�}.`�z�%dml��ks!�c���ѫ�di�'U�lt�E��9�d:1}a�U2cn5���2���7���[Tnԕ�/�!��n���'�ui¾��A=����M�Q�6�O����xʓS�!,�X+:$�@�7�>L�޹Y��Z�v;�6�OU/�_6�A��3Y��>���x��о\�R���'���U�<=>6c��(�}P>!�W��>�ag����5����)�]��K(�����S3�X9R�q�Ն��o2/�z��`ڃq,�/�`�{Q�\E�0����5��\k�ؤ���� z+�$�Rg,R��(ߡ|$24?���**�b���PN�k����s
���$Rp��Y���	�J�FH)+�GGh�IPĤ6��G$)
��,�,�d��g&'n)Kށ�6��-�<%¤��s 3v�(WAσ*������)�s�|+#��]�B�l3`�߶�wI��xލ�o_{���.���u9�hzT��³��Bm��0 �W�{γ8X-�Ղ.�I�:�d�wj9F�,n���'�3W^KF65���g��0T�+����^�s��C}��F�)��˯�i�L�1rͻZ�� �}�=�̔0Ԉ]vn���uw��B� �����u�v����w���*;�ϼ1�w���ڻ����%S`UPM�!�e���y�����31�[_��r���Vs��|=cs�0Dk^������"K��n<W�FjX�����>8�{u������W�[u��6I� �������o��6 (��m[aqL��:�G���H�ĽOl�R��U[�d\��<�[���ג����X릴/��Mw����`ɟ�gް�:��>���K��l�}�ffH ��T����)y,8)] �cu�1t�+��7獙R�ӌ�W���tg������iE��e8d��M�c<6�[�i��B��_��Fi�x���<��U� ���;���0��
���( �62ξ���T���&�b�9u.�6��,�a��j�n	1���;Ń�ݨ��S��S�ZY����(�6����Td&�_�T"I�I�l�	ft���C⇄���2�Z�V��>��Z���<� ����]�������� ��km/z!�c}��`Y�R��S.I2y�D4�|)V�ә�Ac ������mQB��8$d�����q1!����'_O����y�׈��H�����?'�o�P��.�R�z*��f�n�"�jܞ]s�"���g!%��Pt��!��?,�^�=␑y淁"]�f��j-y��0a�}}4zŻ�T���r䃉���s�4,��f"�~	ӷqb�xk���}f-\��PZ Y;��W�=xܥ?ަ��I�K���}�J�����ꭒS��"7�?ȋ���]w7MYZ���%��&�,���Y�'R�C�i������������t�+EV�F�$���t�N�V������~`���UV�����\�.7��P/0]]��	G�HiHm��|	��[և�����E͟��}�c"����(J7Ƹ�5�(���B�Oa�|�����w{@�=�����.v=�-)�L����gZ��a���M�I�N��P�h�dT;�з\J~�@U���(2������	�n�5ʢ[K�����7�,�ڜ!�cDs\���>�qY�(�U�
؄|�̂�uH�Xw�����|�gL�k*�{u��k,w9�("��^�pf��Q���~�i2�R�X���L�j�7[h�v+e�Fz��Ŋ�Y,d#)+�'�O����AL��L�v����Ҁd�QdZ����yxX��"��G\�e�e~aкT�� ��+�(����0�k��BI��<����j0F��e��I<�8���>�21��d.LK���ǁ0��*}ʹ�$��D9���}*г�͑�J&�������~���=�R3Z�}�舩�BY؂�[K|i�Z���IC�#$V���1Z�4���Afun:�>���a�?�W67��/�\OaF��C6
�9��q�+��W��۰ �.��]�¶�X��TCC�_6&��TI�>�Ȟ�tn�����]��F;��tCJy��CǄ��˴�F�(�e �@m��l�ȋ�� ��8��e~G8�Qt�BR�{a��4�SgWj��%Fh�&�����mѬ1O���?�*���{%6:��<���X�h�z��`,w���(\�W~81`'�KM����i�����Y��U�����'<�?��!>MRliW�nO�EBc.g��Y!��ɹ������������)`;QCM�u��q����w�G���⸚�@��T�$���QJ����	�1u�����c~��J��Q�<���$� ����N'��I	�VcZ���{K��>kX��g��CH�E1��k-��sO��+�X���^��=U5��G�	[�.za1��U#�B���"��/5c�����)~�I��.����� Bu	�B��у<�J�9�|�-�u�M�����GS1		Z�A}�R�Y�E��[�u3�+��9'�N�!0:|:������ӎ4�/PQ�:�n�jk���7����bZ���M�G��xC�@����82���S9�2�������7,�)N�^u��H�I���� �dwt���0T�5�>�9��s\�)����5���#�'����; 7}�������(��L�^�����ĉ�Y�rw��h�"7�����@�Lm"ti݋��CU2yK���m�}zS�X�$چ�T=k�F?�zei�1J�=�s3ja�F&�4̘��Q䂐���GZ[��(�h���+fC�b�O��Fx�3�NW�*Q�N�|Y����'66�I��X��w9����CpHfN{#�`Xa+gǃ�`��u0�1������D�ui�K�f<��%��&���p��]��k�3I^�6��t�`��`)>���u�6�mҹ��aMPY��zt�7Z�*��Dd��woF-H�����L�����RT�ϛ𬑰]��Ig���i:���YH�����iCB�J�(q�@̱y����jPtYf����ݚ��C����+�lO���̡����ۿ�ѧ�9Mׯ�Q+����K���ys�%���V&��mEf�l')�6�B҆А��B&�6�!�g�=Q!<L�]��L���/���c���Z�i!o�mc��ܯV���&%��
��x���H�t|�����N���u�b�
�Hmm�`mZ���޲1��i��a���@�6�mx$࡬�7��&�+�}���;��͗N�_n�x��p�$��"�e�
����J��sL!�y�{k��U�kUUv��%Yax�m�%g
T�i��Aٌ�tk�b�����E��l���.CC8�R�(���:�9���X��X#��&�� �(�[����������KO�%����6L�)0}���%M����´;�i����`xJj(J�(F��V,u�/3e�?9)�rV�u*B����T��J�Q�����  |+������s���smSr�?7�"��[Iّ���jي�k��"�|��+�I�P�Z�)g��,m�.=�k����-�j��u�.�٫P�|	���s?��X���L�B�T�ű�4���1���<�'�� /N�[sR8Erж~�����шr�4�eF䦤"k���������{�|���MU%2�����I���X��[���;j���A������t�/e龼�[�滵V/���G��)�K
��4~�[�
��Q���d�H4J�/����ݾ�����P�� 3i�6��{��x`��K0��j$g�ռDȡ"Im�B*�(&9�S�B���-���r�az~�t�XE�g�'O��)�IK]����v���ӛ���(55ҁ*JY��t�H�_��	���7ɕ�,�9�v����r59��������c�>��]�\��8�����զp��*�[{����og�'�W�S�\�zF0�K@E�����w������뎣s���4����=��i|b��76��kkq�#����d{D����s9��K�[FC���9n�W�_n{�*�*�g���.:4Q�'�5�v��ָ�����I�O2f�iE��fY�%�&�j(Kv�3���tۿ��m������[<IZMNk���d��zZ��V4f�9���0~����:Ϊ�K�9Y[z��;[:ט]XqRT��m���ʑ����[H�6	��'���߃���I��(��@����.�ʩ����ĺl��]�n�Q��K�Y4���*�o���ث��i�*n([v����r�-����1XȻ��L�C���Ј��O�deY��l3�_�ӓmb�<>hMF�}׍�U2�}��P��0����\]�2�>���+�SY�!y+]��H�y���p*������ɴ]�
-xX�b�^S�fv����" �]�+n/�G�:�*�M\�&,áC�,�	����	� �̇�<μ��ѥ�&�S����P��k��d9!�(�
�AV�J}SI;c&����'j?X�Q�Sp�	܏a�1���t�И��je7�>�vY�E]��x L�oWL��x��l�X߿�?�����wB���
J�^%�I1��ep�Q�s�m��G<KL�P�|�M���K�u�f��O�n���g�x��u[�W�	�5�|�TZ��!�(�+�w��P�	.f�&ė�Y��L�l����'�PF�jl��*���qa%⣳V=l�ڂ!���u=�����+�s�G�P5�􉼹����0��I�'��U<�|�zEk�OCJ�a�増��)o�rm�����f"��v�fX�Ub�^'G� �z^��H��g�2@��%�@�ɑ�e)�y�}|YN��Ζ�5U�
q��Ǉ��IP��1�9�(�ک@�t�݄�JQ\Έ���f��ָ]��$[~��)�(Fo�b��Z��K6���N�"5��T�'G�=&�,�&�bl��Ļ�p�*z'S4�`�8̈*\؏��N�}qXr�֬[e'<�S�o�--]��&�b���.�w��(��R�L�9̞�r��ॖV����<���d�a��bid��OK}ǻEӽ���R�6�yX�?�^�'I���y��T�3	R/���0g؎��𚮠!���=0�j��>�o�o�o{9���@]T��T�<�&0R��,�>�ɟe���4�|�)��'q� ��0�-�g���-]��(߷6�6��߬���G��0Xn���D1���U�y���֯7� $zӅGn��:x��^3�(��E�9��>Ӫr!k��x�~D�4"�5mk!��	,H�+4I����0�(l'�Q��9�ܷ�2פ��b�����`~�`Qh�/:j�)չO�%p��g�c�z���M��z�}�<�ak�B����q����n�a�:\#�<�.���>#T������*Y�Y�w�l�I��$q��D��ߑH�6Q>����|%xZ�C.a�jh�b(��-`\���ߟ�WiQvfZ"#�v˵�l�)7����g��ʏ���l4T��Ծ����{��� �zpܘX0"9H���7�V6�B����$z\��$�+e6B$|�����3Fu��Ix�ֹ?'Zg0r��>�}� ���z����/���	ȔP�)�����Nd�ҋ��h�a���E�3թ��<Ry8Ӿ!V�����c`�>1�P� @�%&Dͦ��ݳ����.�=[ޯ1ag�ci����F�F�w/�ǘ�@��������	�z�m�uv�S����vr�zE�Ț�$N��� �8K ��E��lpFJ�o��VTk=$;����U*��I���ND�;^�u��C�K�+��㌣{�`�li9~\���m�������h3D�G�c����'��K�j�4�yn�+A0�7�,����M����w8�Q��|G)��kl3�@$��*��pX���Q;Q�p-T��P^!���U:��^��N�W�?��+V,��ɛ�~w�r��S�׊���H)Ws�B3�^L����Í��C+�'�`��5�p�wu��%3�~�Q��tn�^��3qs��_F�����;�c�p�����!�uɊZ�����^���{��҇����%����O���C�'�%1`��J|�2	D���OFǥ�ˇ�I+�����p����2�o��>�B�[��_i�VFnRZ̼�	w�v<���Dz����#��oR3C��܈NG��Kq���ΰ�S3��f��q�I:d�-���ֆ3D�'�C��t��i�>k��_A:Peq{:o-�HFG����r�g��tt���:=�!� 6 ��p�43d���IX��֙�9{�
��#ߛtS,m���y}�����LϪ�f�Q��D�v}84P>JՏ�iuJ�u����Mfr�9|�f�&��E�yӸjd�F�<�B��U	$ڥVvU���Ww����->(�J�k��>��s��2��D�C^�W�7�g�p�|����f����];j���*��&�s�"��?!��g�G/�ѭGu��`�ྖ:���g!:2�d"��8 G������)^T_�ݿ?*�������4@��̒矄�'�s*�RB�;n�$`��e}r����Z{?��ʣ�D�i	�{�8�؊�ʅ6IbI�%��s�2�t�d+AOfD�se \Q^T>��臋����痲�2��H-}����N~s-�������,`�`Uxd_��E��Փ�D��4�a��NZ�'B�ɝ�j�� �Ǘ@��R��'�CYZ �����|�SUo����W	7�ض�6sw�J��Ǣp��Rb���R��5��w��}!j��u2��n\��_ҋ@��z��Ϟ�}8	��P�@�nr�A4=�8.��~=�Qg��_�wGֽ�R�B����˝�	�
F�3�f�d��llM��.�f���
)_�Om����ih`r��ܖ�!G��t�!K&;��j�
i�˭�;d�	�1���8���L���*����1��h|�ֹ2Q0ï�ʄ[3��I�m�����<T��-1�T�f�jn��'��=�`p"O�t~�B�)��+h�����`du�����n�4���E��
)��y�,��> X���f��RMh׆�_�MY����po��"C�LG�M*"�Ilk/?�$("k���[S��g9�M١��n(K���٪Z};Dm�c���-|��mL�<���),�3k	��M�\ws�>g��[�,H�ʨ��Z:$]���l��ɛhf���fy�r�d�_u
ʁh�/	1��XN��\���gƛ���'9�j~i�����C;'',���y&�C��Ȭ�*쿳��|$�ӑ�� !.M)|�,z������xCԸCR�tS�=94��߷�?N���%~6��ӎ�f�q:�_���}������6��R��^�n#���T +�[��1a�* B��n�zSw��C~�l2λќAn��,�@{�6\���i��;�tg݆'���y����)R}'�g�|�淌j�ٱ2M����2�N4I3
���2Wڋ�{�}T��Y�m���7z�B�#�랗�(b��[���K�^�W����sþA���sk���*�ng�C[[-���.c��B6��z�=6���0���@�`f�<��ld'CO	N��R-ÂS���@��֮����"�R6/��;�GJ��쭙�$��ﴵ�
L��e��|���b��,F�Z�]�/;v����3/~z�ݵ�o���ޑ?ŮH�k�ۦȳߵ����7��L>sevr�`���ꊡ!�ƫ>����;h���ې[D�&�_�a��gP͗����my�b2�֒?�"��/~�'�,����J�+1�g��fkl��(tG/(?�`�B1�݈�Qp��гWm�N�`|��qP�b��m��6}q����%q3���Ds��+|��e�\�d���*�ߣ�M����Qi+� �Hw�D�J?ka1v
������8&��V����(�һ��<hyiZ�3�w�G�)ʴ��/�$(�~�w>�@bz�q��=���"�����.#���;ʌBV�2X�A�������+ק��I��v�G�U�Z���o\��m�2v��qke� ��ʷ����b�
����e��d��c��Z�
���0�����f����Sc�_����d�1ecUPq�8�%?P������J���oU�2G��>�]nV�	h���^L�<���3poMQ!��� �][ui^\4�D��3�wyy%���<��ʽ��,��f�HRJ�����U�e��������o�w�A�^�x��/��&��f;��p�T#[��\�z�/iϮ&��Ǔ�笤%�X�ҹ!�T�y}.�=J/-F�2�جFs��������4BjQ��c!�S�t��{u<VU�����xr�w�!�2fV����8�P�a�%�;�S�{	����ԁ�(�yT�\�=��*"�EX��0���7����	M�0� ��,�_��>�M��'��`v9�!ύ��Re���-��`�y�O��T8+3�y���[�3ӄv���!h�@��"��`��3s�"�]�Q��0O*=L/��WM����X8[4���GU��-��"'�ϣ5�F�@W'.o;Z,���މ�xkSU龆	�kz����K2ϐ�U�9�x]��Mb�cR}Yb5}�E(�Ũ��K�y�H�L~��'���u��1��:gC�-�+گ�?~ui�ș�[�6�Np���W;2l�u;��+��"��2l'�^����5G�=�o�E�����#��N�s���q�Y�M�'D|,Dvr�N1�SY��#�#j|k��cUޡ�,�l���#]H��߁qɳ��y�����0u�}�Qգ�%���	T�l�
�O�\��w�MD���M��#��p�^{QH�ˋ��io�K�F�f���z���h��w�{)G���Uv�"*�yV��so����&�a|'cK꥗$q�U�[��n��"4Y�^����b���pŞ����� �d��ȠRsE��l�?~zJ�bS!?�q���ʸi�7�³��V������e����x�4,���wlʲ�����Z�k1̣N;���59��mL������B����\����o495}AJ��s���86�����9)�PˉQ1��x+��߷� � ƈ���`�/z��TM�Q?�F�#-�����w�����Ʌ�6vC���7�y��@W�O�ñqZa��dÉ�(��-Mpɹ��w�E>�un$\q�Q�D|��$c�k2Nŕ�����j�Ik���JdC
R��d��[7��Q���b!@`'ZQ�&�n��@K��:O�)�q7;Ya�q(��<]4�%=��l��9�j਩ʢpm����.��!I �IT�B�@z�r,_G�T�o��B^��Q,�Z5л�	��%��P�����5���P �Np����tXe/P��&L�p��eI�'���2�=z�.�tZ���U��*dj"�-�W?��zn��6�T�H]	��̽IG���wZ(�s�)��5�E�=�y6��j_\�p��Z��,�o���Q��<5KBu��^J��)ʌ2
z?E'��*�`\��Y�9͜�ݡ�����{��%aV�Q�������u�W�S{a}Y#N��(�c߻����9Sh�Ww|��p	b�$|&%Ѹ��e#C9d֠�΀[O.v��}]�r���ʬ�����!��A��5v[m��ٷ��x�X�����#�9�� ~�2nI8WL2��.d�u`�$��tէpu��M k�a"��m�8l��V��BH��:���W��E�j}��3�{�������e��ceKL�`-�g12Avid�y� zuA��lv�K^�#ΉZe�y��ՙܝ�R�瘦�!dL��C��"���=�/]�w�-
��Z�VTt��F�։�M;���0n��p���5�	dq`�p������x��M��.s���Q�N�;��B�s�����C�g ��4�ي9�>O,�U�:W-����jd��'*}���;�",S�c�����D2��փ���"7)��~���
77�#�׬��@֓�|���;�<��<aӚ\�n^��uR��o& 4��Upr0��g�X�i2a��&��5�9�ڲ�f���~�i,!s��Pj ���J�����K��qk`�]�w�)�(6�����Tn�DY�h�R�Z
zۑ�5"Q�u��=Ҕ��-}`��Oz8��cM8Mn���k!��=K�<�W�s�"���I~�a��=ʹ����A�d ��{-�MQӬCe*v��q��y��M� �"%S��mF��܉�LZ��ti;�S�3�u�LkA{�+�-��7L�\��*6y!rW������=a��i���E�(�<�
$���ѕ�[n�f�'y��������<���3�g0^����~���#u8\+�{�4C(b�w��j��$���P<<'�"<h���n+ 'A���i�� ������Pʫ�[=K��m�9\4��t��u�0A��*?H���������ԇ�[����NY��@!���L��T��:��C�|�6U��.��;P煌�2&�y��������������j���t�If�q0�^u�o�A�E���{�sA��I#xLޜE����YX�I*ڪ�-��7��}�� ���j@�)�8���7�#6�����g���G� �[l�&�u�[��C��������Wv��bf��L����+�̖��4�{<�ӏlS��on�άXP`���2��^Pȩ���(7>n��m�)�5���ja��Z>���XKY�G]�lܴ���h��u�1���t7s�u��1� �r����r)u��3;J�aW��:��+ں?���S�_cBFĴÛ���>�����:,��������.���,���@*��uoBn�7#��|�����f3x$<@+�wь�j���z�`��6�6�dGwBJs�W3Nm�:�B���({��#�`�?- d�о�۫ �?�2)�f�8�Ρ@����R�o"H�MM9��+f�O�/}�N�_�9�%f�����;�@S�i�k�.�xזr˶w��U�����3���r�q� �2�������.^�	$����cN��ޓu���X58%�D0n_ l_����	n4@<|Y� ����Z[q�n�Q��\�h��iHI���.��ϗ����4�ʦ2��.8��x�]sv�g��	���d�)I����U1ϰ�at��m#�7C�b'z�*Ɏ�ꨊ<s4ց���TJ�C����5r��eN(��,��~?%���d���o��X*�<�w�$�[M�*���g�g�č�G���a467�n|�M�!����h�[]-��}$���R��ًD�$"���2�~��;�Y-vvLbn��\���܁$�.�>_/��J�:B�@�i��� :|�%��L��&|!t���6�%��,�Ev^�{�a��R2F
�:`qK$r~de��,�m��F*��	�$�}��F�S��5o���; 5�1�?M���C*����@k<3�r�@�ұǛ~�Qv{�� $��5�{3��E� :�9g0��=�So�N��2�)�|0��\�����x�L�ġT%�!��@���9�v�j������0*Ѕ�iOt%{���kX��!�G<XK�y��d�^p��b���J�{�s��Y�/q+��n�1��`ޣ֝�ɟ/7{D4d���%�j�\��a/��]��LB�>Dg�O��E��-���Ϲ�"#�nx���\������ᢺ��N��C��ݹvȩ��������X�7�AS�V�^b��&qGOh��R�0��%��?���b�ڷ�(�����݂y\�p��a��������K�j��l�n��9���,��JP�K�>�|��F�J�M�Z3��(\����j�R���7��ؔ'J�����y��G�^猟Ừ����\���p����˫Ƈ@�X�F+�6�0���4����U�~��e�-��(��-�BiJ'�ً�6���d�QG�'�ִ��W�Y�������js�V~�