��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����xLM�����`,5?p�"���N��}߳�^'��v�Y|'�XR��f����mM�x�p�xV#ڇ��76{��)����L���h�:��+A���9ߨ-� rā�SZ )����C.��&0C]�-��[�3�-���+��պݣ�k�J�vo`�A�����f����u�X���v�=�а���]Q�Wۿ�߸�=_Q�X����j>��Zw�K��SvX��ƥ.���#�����Z�0���#7{��\S$��@1I�QX~TQ�E��db����۰� ���>0�%�9�j汈��}��1� ��2���h�G��SeY�a���	'<x�p��k�H`�H�j^y�0�s�78+���ֳ�`�R3dW��_��{p[�?$�s0��#�zS�_��bH
�c�p�IL7]� |����Q�� ��Rr���=��E즕2%�����`�^��l�q-�]�p��jf��Ӽ-f%H���ȳ�>��+���M�71��4_�) 3�46h�rb�J�W� k�h~K0�>P$�_n)���5�r�j��W�J&޴o��$>��6��ŀ�;A~<6P��K�~��f��*I
�Z��}`q���ApC��n���g���3��-�іrO�mF���,�$��@�BI�q�}��Ȥ֐����î�䂧��@������U���vU������ �T#K@f�㯁����|95<@���+�-�)�����K���FI�k���*@�m&���
���ma1[�2�u�I�\�U�yu���o�|��2����;�W�W�}P�K>%5�'�8���׫=����k��,�t�M�0�8]q3���N���GvZ�i�+ C�e
��Ќ�S�v<%���q��e_��
�k�夞��>ZO7E~��5k�TW Aod��eE���G���ɑ-'���?�G$����ќ����8ɸ+ 5ʗ���l�d��,�J�
�^�3b,�����J����#n�zK����z�&��;|�\�^���'e�W�����">�w*	FO�Δ��v�ƺ����U˲L�[f�$*�f���}��6�T�
�/C�)�]|���A|b�s6�v3��O�2x�-W	�����	D��5A�e�����[��Z�o��R@�eԁ4_3��+k�%|FARG�M8q����d�˂(���U�on���d0Ͷ��"-.�i}��t^�!�}E?{j�~@U���{�d�b:��<�XF��U��T;�NW��^q(k�s�1#��p�2ߖ8R�c�6]���鮶��;������� ��K�S�o^oFjDբ��o�Ct[�}�U�� ���B��M0}�F:����޳����Y�)����,���Ǣ]���^f�6P�ť�;�jɎ6)�����m�:8��}Z��4ߧ^�J�tk�hks����Ig4��T���A������)����y/|u��g~Y{��s6Ba��Hԉҭ�b+�HS_��w�Ch�H϶Q��S��F`�Z���r�H���B�4ER��II6z�q{5[������~a%[����6��4����3r���]TIc�{*(t�|DI!=�Z�|=Sg*홐�W��bd�ш���^H��]L}3}�B�0�̷{m�qn4���?q�Gg!6� �[O���ŋ�����������{�󍴦��Z�f������t��[@ܣ�7�H?��{���,�~�w�O�,���Arr�P�,�X��s�g$xY�*UO��V|!����V�W������� -I�%Ms�l�Z}F����1��ם��8$����P � c��Il�pʪ�Yr_�z�E`��U�����XM���Iv�B�#�ɘA�&etPKaY��y�V�1�����G|zs����X]��x�(;y���� Mp�O
���;"���ڜ����U��i�Kix=YC��ԓg�Ő�~NU�cj�)����Yko���!\���F������b7X�ф=�!�Tb���l�'v���e����;��.�>����Q��}}(� :�q;��	JDq��=ݖw��T(	o�`˫�	�ibΦ�k��֐l��4bR�/D���i�ȉ���'�/(v����ك6y�����.�%9R'}T��(�]1Y1b�}c�ۼ�K��s�|�Ci�8�j��R�6�^��\��.N}��@WA(�&�o��@�/���>i
 �j��5� a/����v��Ǌ/����a6�sn���5�q����/U�c5��[7s1M��y7V�P�3]��G�l�W�{Ny�@#�ђ(�E�����Fc���_�&�&��Yᮟ^0��g���KG�����3���u����A��W��)��ؾ� {W_$��3�"�n����2o�rꇒ��1.��i�Ru����\��R��o�摅fN&R�QS��p���]���VA��,G�o{�M/4�+L��fx_��<l�rO3b|�l�x̗�?��)0o��{7/[`�1�w>�5���Mz������9�3�#���F��\ ;@Ywѻx�ra��lkv �9��F���~������P� �tz�綘Sb��PUX�?�&W��e�]����?e��'������7TPx��BCrM�k~>���ڤ�N��	w�>��uu��D����*:����XU�Ϲ9�+�U<�����n�0e`�=�$'�'�%�2��r(�<1Jƃ�u�b��]�?�Pa�����쾯��\���a�ϙ���Z;�<�D r�е��Fm�f��V�(	O�2�WF��$Y�L�y�U̿��d�5S샪���$##AJ_��Kݻ��ͦ�4���
. ~E����y���)�[��O�С�gQ�Ҡ�$��Ad�)E�,�h�ر����ma4SEm�b��!��d��KB^���B�e/�dPB��#9&���ȭJ&[��$ݚF	�2�7U�9*�)�#��A�2�^aL�:�bCE	Rq2�Ad'!�����;L�v7�b��\�WDjq�p>�Tf��1(��3�v2�){Lp�l�e�.��������$\�o��s+�fq;�n��[�a�[�q��� �E������g�'$��檝T�O���g� �Xaf5k+f'�*����2���)p�KŚ����B�眻�2|�5�"nKi�QdQ�~p��.�t��q��xQ����ie�ȁ�o(����O-��&bm���,g�9��Z�p���D3�k����"���V9��ns��R�X����s&wn߼�RH��M9҃�'|�8w�8~3���;ލ5�*c;ͯ����:�ֲJ�A���*��)
>�6���T��l8;�{pH����Ί�9:���� �2^�5.`ꨓ��yX�Z��JJr
�a��_w�Yy0��0�)���(Kz,U2k������5 �8BH��a[��[��V����O���4!2��҆�AI�K\�U�2L��]y0r�*A�d�����͉%��!OG�#�BC�L��V�?�*ڱ'�X.��UI1���8�����!��%���<�_R�S���?� ��o��}�L���hj���e��b�4��0+��H�HX��I���f�r����g�HL�qw�[���+�p*��C���g�4�֧$&D��
����
Wc?��,��͆/~A�j_^@��oJ`����Xb�gۦ��G��h4mt�;���ꢘ�C��`����""Nz��}UN���"k��߯����(̃QN�t�����ky�c���6;���E0O��W�a�Ò�R�s���[l��u)���I�2{m	��с9�k��]��X��;&�T	2~-]�qF,�,K<����?1M����: R�b1��X��w6󆗮�6���L_�Sp����]P�^\?���*����j�E�S0^*�C�z0DLj�"���]�_my��C�h�E��Sq������4�qr���ڳw<�JEm��^��A	��mA?�����5�3b��qGoY�wnP�ǒ#�]Xŭoc��B���!�*+�=u�kM���ߘ��U�J�hB�����5�\9ʹ��&�i��â!�fiw�ͣ��	�/;rg�N�E	�C��o��'�'�#w(E��m[���K�[���x9o䣐�;S=N̴���.��)
6ٯ��f�e��s�~*3���Wu�������n�K$�7v乂p�ɠu����q,� ��7�A�)/�P���=J��.~�u�-�7(����ɆD3�J�:���A������#�d4i]���4p��ad1�RR�Q���j��ќb��Ʀ7 ^ӦއhW��O��-W�I�\4}�u��&�l�g���b�p�Q��Մ49 4�����c`wM5�э�;&���@�r�n�%�[4�H��`@"g
^i%����w
�H�N����n�Z���S��g�d�H���B�-o������eC�)��1��PWL$�;
�&����OGx�>������+`�'�r4vٽ�����?�Υ�n���v^^<�t7L#!�dؠU��������}��_�@O��d��K�U��C�d3�{Ȁ����]Za�4��n7�@� ��T�θG"������7yw���-_�[�� ��x�D3�KV+e�o�Ì��/�q�ɊI��t4��'�v��+��@6_��JO�l^Ӊ��>�(�&
w\m��/�y�&��wH��/�k�M7��)�$M&�;F�n	K�/��W>�f��hQ�~�6�t�����ؔN�q��Yߪ�;��G(���Id�����3���֥�?�6�?�b���¦������|�_g�ᛊ�^�ۼ�����ߗiy�n�v��[���vU_	k���]�Y����0���^���+����$��ܣ����u-��a�㣩�4������
8�p��	�K�9�я�STg�f<RQBM>��c~�'���lo,��6�{ވ�4FʄB���YU�x�a�c����gn_nť;����Ǌuv�R��NS�<f�|�{�����(�
wy�^迠P���0�~���G�m���A.5���KE㄃�� <���� TNh�1��B���F&[>���~C�$�0��Gu�6&�C��o]�%���R�(�U���5+V���̗	��%��p���8�>	~������jc�d��1�9��ݩ�%�%�'.M�<����mb3������-S��Rk�Ӡ�3��������Y!�p�.��)��@V��`�#^��&�c�H[�O+�`��06��r������v&�=�3���ؼU��J���j��1�|��*�
D�ƋL�kᩂ����%B��(�fn$3xqtE�\e�t~ �����7��Q�M=:2��%M��h )�ÜJkc�3��������z���(��/L%��J��j��0��9w��u&���� n��r�����-������w��E&��?�  8��4��o���>��,�z�[�a��p�	:����Dyg��F���,l���I{���kIi�T��;�F��q��-��0�:B���">�"�V�R�����~+8l��;��,�[��eʲ�������o�������9�ѻ�+�q۾�`�n��#��J��f9и@��A�s<,yZ����h}nT�Rׄ�>�\i��x_].����
'��j{mL!r��W�dW��G�B/��0lb�U!~f%-Q���~ �9��H�A�$�������n���D�-�ޝ%�b����.{8ӎ�%@ѹî8��}���ٿ	�ρ�]�T;2��a�0�8�U������pV����c�a�<$eO	��n(3���s��i���#Pr��o��QHP�n!�Ử�4d�P�Qh�i���d��-����;�I�m��h���GZҩ��g�?ZT���Y\kF�#��^1���"�����]�	��#�յ��2�:�m�$ux,��6�uLԷE�(�%���׬E��B�;�2�t(��5�ȡ�̕�����Ogr��c2��U��̉��U�\�b�!P�d����hhٶd�����.���N]E���s��k[QՁVRX�"Z�~)̥���Y��{���%�ҎO���>_����t��q0���Ap�&)�_�z�
~����F�6:��o����>�Kf���Y+��1d�;�&:�܇�����i���	��f�eM

��t	�Vg�0	lzq�}|4mKr�l�Ǉf����͑�G���t�os	~G����h�_���_���Ջ��fh< �{8�Ny!���p�����TDy�&hZ�=��� �mF��?
��z�%Wmm�v̹+`A�u����}8瑋��GeLnc�������Mr5�Fw�������*Nr���e���Ѱ�u���_��ĉ�������H\�২�w���*n�d2␠{3<�|�b)����?�D<�k��J����z5�G���(��y����x������:������N:���,fb��S�~����+ln�}V޸�GJ�Nq�~���?ۚ�2۲�
���`��?8�:-��ϣ��#�a��I5}~�^mb��P*�PlؽTk-Prn�fw�*F�^�Vy&@��\_I~�_d���H��f\nùH~�7R�\�0��gBu�͙<71��������u���Ǎ V��;�r��6f��Ʒ~Y.���l�;�����6BҷE�ۖY"ؕ[�X����3����<�ij�q���4	�W���o�4��sCX*O��b�[�5�+����] �F���T(�J�����``�&k��b�HWs��5�K��j`������_��6��ׅ�"����L���w���������=%���T�����*��.��r���b�u6��:�st�p��C�N�XD�@�k-��l�f��3^��3+a
�=�̱������x�3S�nߎ 	�Q��,��xSi�v�:�W�D���ǭ�M}���,�!�M�xhJ�g՛���������-)`k��_�=Vc���D��ƨ+��AY�s�|,2=�v�	���WA�IN�� �f&*e+�,�������3a�D�L�L�{�j���L��x��F���4"�̃��45��ӔL\4�=s%�E훭���ͺ-����1�ڸ?�D��S]T�b��_�
UL�nv �֍3���{\z6��-�n��Y��&|��5��<�M�z�ݹ2�_���U�kDfނ�-S��S����A�Wt�]<��q7;M��Gߕ�	�������-��L_��*`NU�� �¤f�7�&�t�zPU���	9��
�3��X���!�c�k�y}a�H��Ӡ*l�+X�@��?_A�0�LT���$ �e4Y�Ͻ.8j/Z��vTΩ����4��2��A�LZ�Z�'wo�Z=�������tk�ӇK/��ªM?���&Ň�nG�;���ۄE��������p�E��-�#Z�ԙ�YJI�� ��d�	4&3��oܺi KKf���t�"1_�&(2����A&�[�Na��[c��/n� �Bp&5�}�k�fH~���^7�:N;�������{�{
�S�K���ׇ��vU����c��;Kj:���j�iwt�N4��`����7�ֈ�T�U�H�)�c�9t�`����6y�8����֦�z�T:��	��'OBΒ"�/lh�pb4a��2ӻ�y���`�ޣ�]�F�I�V�r(�iVRJ)�f���6
s���jn*7�����)�Zǧ��.zן����%>��@k�T�1�4�q:��J\ZA ޜ�+���Î�A�jE�7#n8�{�AV*�i��bH����>Rf0�<��L�Gδ�2�֮rG��6��U\���[�����3;J��S�	���ˋ雟4�A�az)Cq^��;��6i��~�n�EV��5���z��ɑ��jq�f0����4,*���W64�g�����eH�Op���	�⅙�4��}�1ˀ�� �T�\�Wt��sgR�m念 �Z ��H�#0�8cՑl���|&	�8� ��Ɣ����vA��a�5 �1F�O��n�/�_K��P��yB�����I������.�/�	���)7Ȁ8�l$��Z��F�F��� �Y�d��Zv�a�M柞Kc 	x3
G)�	�x�zM�S(��[��Ŝ2��l}�
*�uOjS���C¿2�Q9mĄ��^��${&�@|8�b+��=���a���������,4��˓�k4�e����DKr�t��2J��
��I,>�-W]+�@�+nK��^Y2=��t��S��ž�����kHS����/?��3M}���*_�Կu�(�T�?����z��ID��C��ޓ���Pkar���w�P�����OE�&*���'�H-ِ����3cZꟚ75O�B���f2"���r�s(�9~rMw�Ě��d�a�3��2��,6BU#�J�^Q�Y
�ڭ�s�j�ËFf4�����_�VE�ټ��m����������I���fBY-���J �\�|֑7r��g�)*/&7�����6c+�������b$� ��2�`y�0L%�aAA��o�e��lq^;���������A�ișnFV�E̿.q����(�g|l<\Ab����f�V()�3
4�?$�N��򁕟�<T�nL��xj[�c�8�c7�f,
$�3k8�1�P=���6�_��2 �J=k��d�v�o#�}`�����]�1�7�&�U��ORڀ�W�{��V�h�]��R	���	�ͧ	?l�
$BXAE��� ���C\x���]��k	7�;�l�Vk
i�?1���L(��K�T#	)�pF.��iV���dl�U�W	�����-�����p�_saBŒ��ob�T ��c�0;�@�b��w^ڎ�?��Œ&�Kv�%5ʕ}���r��MY`�"�.�w{��?���P7�����a2ZGq�d��8�I
v�����`h=��G�����w��ī�jm�{-U=�jm���_��	����Ȯ�^C���Ԛ���p= ��j�ruAf-����t3W��������{��
�5i\��T�cB{M� ���Ԯ� ���v�>!v�4_�.���"�l��S�&D%�`l�k�u�D�Z�T#��%8��jq��%�4�w���wh���8���5b��5��$L�����a@�t�¥?��bȇָIl���f�W��^�l���,�l��ԳU�Ho�[i[o9���rQa���w��K��o;x\!*�2#����n�Ӱ��c�"�Sj��K:M���/�yoض�7��M�A���y���T��
���%��eG�4���徑�F�s���2�5�k��4���m`RL%V�ϯ��^V��_�$&��B��U&� �B�ZƖq�l� wB��"j�!+r�8�����lajƅ6I�.�ׯ�;rn�o2	n3@~�u�� ����Fzf��p���TT p�����>y��D���y��ȼ��c>ֿ����*_���ȥ�`.��w�ꨠ��т��/[�Ij/@���"  �O贄=ƝeB�(�������,̰��8H�<� �d������t�A99�lNĪ��x�[�����b�	���䂂�=�lk���;Ռ[[h�N�}IA��_5��WJA
N47 �[�`l}�����%P=x����DO*g8�?l�(3�V�`����0!rT/a+ķ��Qp-��ZȚGQ���q�X�*E3�T���8�E�&i�?X�l�^	d��w�Ï��b�n��^�]��IO��Bxʨ��!��S-�J��X<��@5���n�\ճx���,�3q����w��~V�NY׊?����U6*�쫕Эz����h3��n���2. �}D�!���6��v��Г��N�舜��|MjU��<_�@���-3|�F	p�-�P�;�P�|&�����sԂ��e��^��%�a
B��!����a Y��G���l�q�;�cvpf�.wX����Y'�Ti��+�?�"�wtM `���^$��00��,�q�c��:�x�^t8�}+�,�6�qP��Xޛw�/;�Z��)�����Ҽ�@���8C���f*��L�B�gTd������p��G�0���bQ1���HN_���˔bT�ޱ���:�a��F�p_��54,����zT����li��Ӈ9�fFB�ig<䳲�.8�F��g�7�>#=vl��_��=É����*kݘ.�О��<d�|x?�VHHsڼ��|6\`�Bئ����G�j�u)�E���T.m*����H0!Nգ�����>��:�&ɦ��h)���;N9�l$5�Ki�t���	T)|�������)��À��%��}�"��pe���j��j�ev�"��|C����P�^/Zxq�A]
���dܾ���	O�sEȞQ���Q��� �7��8=�Jo���f���6�䳦�}$�Z�|ѵR�����B�1�ef�#���!P�е1w�u��s��W�\6�W��{�k��Ѫ���3�N.���qz�ڙ)�ճ��q���>��؈Z���(��-E���E������]�LT9<m��j)����歫��Β4ئv���lKM.�����i�D�$�����쫣�=�=Ҥ̄�l�y�#�*ϓF�F|��A	s� �>�(/�N �]��lW��PG�:^M�C$ؓ�$���7o��0R#Y/��D`���I�>{�e�Z�m��
vz+����是Z�a�[*;�E_��Li�W��։�K[`"<ߟ�U���1M@�PҼ��^%ۂ�\��(w�8p�-���<���w0�	pi]����U��f�O��4ɜN��f��_�ͮcQr`�L�g�@2Ͷ'���՞x�y[X� �,��D5�`�ƭk��2<]��E^���h�pݕy��.�*���i�ɀ��DA��<LU7}�b��}C�,�}�I嗓FMg���9�
A&Α���m�#=K��s<?��Ip�Qi���Vp���$xr՜�g�I�;2r��Li�m�����j����z���>q�l�����%��\ZG-�ގp�*�� ���7��B��)�����8�����3H��M�N�r��!0�����g��G�G�h��u;E|F������3�@`^�g�l���^Q�׻��n"���@z���$9lj
l2��"�������t�պg�	�����7g��)ZP��4�,�� +�M�4PbV��+*�V�(� �ZfƠ��ZPZ��~�
��	*GA_��#�i� ��E�7���,g��xy���!v�2�O��[
׃3b�z�g?rQ�������z�J�E��:��2�_#���x��r��j�t�*:ūFJIɔ~-�����Ҕ�hcȈ%���������E�`���L+�C�M��,J�{5%���e��\���޴�j+�#��^��j�YdX}\P�]]��zY	_0�M��(5�oF
(��i=�ծ�zÚ��z賋b�ɜ���iaE�y�{���}؃�� 4�~�Ϛ�~U�m�%�?3�
�h���{ed�E(S��a�r񇋧�&6e-��h���yK`�l����9�}K&(^v#� 3|�8�|+��.n�U�]�J���'�?םo�����>��|l��/��$h�[���;*B�T��;�fl'=�쳠Yb�w?�wy��.P�z��v��͡^���<G��,lh��d�-0�7[��e�܅Y/ �d\�D�k���D7E��)w�}�;o � W����i��
�L7l`�ҏL���m'�Q���Ve'in���s1�6F|B@Y��k�p  ��-�%Gb"L�
h���gaO�%�� �30h^�{ɋՑ������O�:FK��UB@�I�ٰT`��n'ѽ�A�Nb�Ԛ��cH�R��u��w���BٽR��C��h�+ǀ����F��==�y�)q�x-Y�`�/6{��F�\x~W֣�W��U��͑MO��Î0��V뤵lNq?�4�ɴ9�pr:>�5o�K�'�$�FE��N1A�t0��21�[�px+K�$��w��Mة�A&�x���˰�5`	 ��Xƃ�q�ݯ�`]�N8!������逅�G|�G�����E��1G>�f����!Q��q ���D����{C�D���r6��0����b��e��ʧ�	Y`c�\m��d	�8��`���:����dU��b�u~�<<�1�d4�����q�6aD!�UO�ua�8�iO�v�
���6>F�ހ�A6Q�Ei�0m[�-<*��s�^�R�k1����I_�DhP.W41����b���n��!��<�Ǿƌ�G�ͦ%�ߎ��b��j�<2���sU�+��֎������^|���/!�.v	���JIj��'2�8Qx�bK�6q	 ri;��X]��h<Em}�������>1�4�;�٦��2��X$%?�눅��[�}�	&Б"��^�����H�l
�\��բ����|N4s�lκ�^g$`��]a!w�7r�|���6I�A�}���N�c��`���A�
��fx��V���,x�YDM?a��,_YME1��o�����͔ѐ�fT��@k�XK�m�C��Kg�կ,"Dr�t�sB֥��b�l��H�V�xCZf��3r�H<?�j.���S��W�㕙��;b�\5��5S &؊�F탖��Y�D_�S|�/�
�Ok~.Z��H|u�&��K���'�G�s۟
v��l	G�΅�X��t��4N�9����`�}�l�\bZ�
T!]�dH��X�=�rd�>S��r��S��	�F��ދ�*^�b�]3�k�Ꟶ��<�(���� 
 깷���"`@鲃�k���<��7��2��Ғ��#����N '�D�;�:pۣ�Q�$0�]���v$[���/�j�������������������-��8՛3r�3�4�~n������� %���+<����R9�c���������y��+�5�  .��Uԯ4f��殡%K��z)O5�����_�4F�\Fq�_���0F�,����_gn���P�8g1��M�{m^ʎB9����fz��Ov+��3-fm�jFRxU7�b���^3��`���6���5�q@��+b����GJhz��f�
�j$��]]��8?R��%��/�w�j���ߠdu8�������W�Hy|���''ﶵԮ��Di5q�eoj�:|7x��&Â �H�oT:��0�x�0-���I�Ѧ,U�� Nb�0�	�!�e����ǰ�����~�Z����m1~�®�:S	�p��^�3l<W�Y(F1(� �9������ �$ֱ;���N��� ��M�FҊf$iEA�q���p���*����R<�����n�T�N�o=8��Rס���Jp�cad���ϓ��V����tݠ��cI�`d� �1*��$�
���`�'���{~�Q�
�0��>-�s�Ń��@�i�ף���f[v�S49h$,�$e;���&S�Z�k���3�A6��tvu ��Rꁳ8��ę��b><t�W�>�~�e�B�<M���nM� �c��[��xI��]����	�ߵ����曭�����esX��Ie|us�m�����r�A��܀_z��C���S��6�����AE�b�4�s��^�ɩu>�(���Wc��6�A��X%�Ò�Ԣ�\:NX�3Ϳ0R��s�A��T`�)s��=�<0;����9u1�F6��`�#Oֿ4)�ؙ=��d�p�����4��e��musq"��� Y�9U�����k�`e���/2�2�s�&�IF�G�s�r���}
�Q'5�AE��*�A�S���lZ�%��go~n� ��U�"�eA������9[�|A�Rų�ur�T�Q�O�� ?	��w�K�e�;o�u� �q�*/`x����֚���M�.@��ǰ%G���gM�M�w�mF��΂'!�y��,@8��(����4���v�.:-j�}7�5' N���� �SY��L��!���C��E���T���;L�?��h���إ��zߩ�Y��Щ��\�]�
j��wI����*� �F	�	�5m��޵@�%֛��^���������>�E��
R��(���e8\���N�k��h�X_]/��\�;�_�塶	�GOg��l�,b ` �XccN.�M=��y@PŐ�~)e�ĕ����Ġ-�I����,��?oϋO ��s���������FX��Ri�}����軆��o�6�w�%m2�_i�`���T�7��p��Ow?%4O
���Hu�[(%����gu01[n�Cd������h��.�=���2 ����z�-��{�nO0�ZW��=2��OC��+��&��B2 %I��
7�.��;_k��֣~����w�p�~�5�Gn�C��j1�i�[�zC韡s���r���.��m�@<�N�w�*
�:�ɫ~��-��/	B{�HH�I�iu�ę�[}���n"i�r�+� ��%����yG����ϡdӠ��􍱯�PY���NSN�3T�e�t�����+��������܅Z�y���.\��+�K���������`G���R�!�LӰ
��9�@����s>M�{�Y��)��^��n�+�${_�a�*��p�O�ɷ(�@82j1m��VI�j�E�&�.`93�R�a�w��AK+gގ�cZ����.�ڽM!,���������L��M�f:�����s�"Ө�Q����4�y)�(8�����2k��{�dG�ݱ\�o�3����ay0acj3�ȺPCm�[�7��=� D BxS�U�拝tWݲ�Ma���D~�[�`���%���irm�Y�ggD)5 Rb�?j,��ZT�F$��W�z��>���O�0�b?����?���J.Ǌ#Q�٨��]Xw������wk�-��w��'3�������.�s����D-�rq	�`��(�����qw\�=0�q��ʻd��<�^:Ɲ ��hg=����m��
ȸL��T�m���㋻jm�����.��-�[c*�8@:k?m]5��T'e	V��o3;Ș}@�"�(k^����������!̀�itu$dOEJ��Z�������X{��.�pk-�̓�y�
��Z@�j�O��2������)J3h�R�Ś�6*�`%�.lQ�F!��D�X���Hn��Q�
Wn
K�Kc�t����	QQ�@���sj%&΋�t�X�{�޴Zf�
���qVU��0�8�.�mڇЏ�w�R�r�����>�k=�7���p�WZ�Z͛F��(��m�,��ڣH�_�o�U����V,��n�;��G��o���7-�mBEwE<Q}����5��;�{k5�h';f���fl�S2׷F�Mh����*G��P����{ԃ
���� ��KB�feQ���(`ܦ��S���H��o�����N��K�\��O��rV�������'$�>���e:s֨'+��U��
O?^r?������ж��-��<$�Y��1ӚJ,���
;�S�@L�����<A{w��M��u-�u��Z���[�$�\�O�����s_Mȑ�X��d�13ܕ뺟DP��q=�i6�B>E��^��L��L�>d��8�f���m�&L�z�>�����-v�b�2RG��,�`%���[�:V���8��t�2�,���a�;9%�������{er�`Id�(=�`���>O`��0x��l�1�;nmt{s��-�sRs��:��qi�p�[�jd�.��ǂ�0�T��|��b�5U���
; ���"�#��+��K���r�Y��/�������,w�l�w�×��Fݜ]�#d��l{���2<���q�>TOmW�>�) �jE�>�|��G��Z��ݱ8��^"�mos�#*_��)<r�QZod0�$�n��WS$�w(a_��8�@��%��4�6<x>c̿�c�&C�X�ԌV��trտ̥��rCe�V�cQo��<&�%������E��D�Рz���o�"�*��3LZ��ם�c|&S�[0�V�P��Jo��ʱ	���5�+��<��R��xC6���ux��#'���gU�4���/2y��$�8JH���;&5"�64J�.��<͟�v\e��5��S��p󪐸]��o<��|	#*��t��yk��ĭ�N��VF:�f��͝�_��>�Q�_��	᪫١�&ȧ�t���>R��^��s$�Gl�>?��M=�`��}�7#���<�84G��1��mU��N+��w�<�D�}P�E��`��*�[�Ѣ�=*�v�u�%z��]��C0�_Rġޟc��'n�#��S��P�=�L�{>#?Cc1�vh�I��o��;�*������7��Rb��@]]w	����Ө2\�)�Д�5�p�L�1
b�ڜ*��7{�� 0p�w�t\b%F�����^^��d��?��ۅ��G���My�i����ӕB�J��P:ǐ6<�?R���*���{ڑ�b�swj�D���k�Iڪm	@	I���|qt]�u���Hr'?H������o��C��>��ǖ �bV��qUs������	R�7�#�w2Z�M�m��_���	�is�������]�)��"�z=�p���7�QM�6J!�n)�����wjD�
����O�:}hf��@���⸹��$����$�|�8&�)�Z�@R/�*��H�J�K���e��Y�I�BϮuI;�������m)��(�<�֧��6O]>G(�mp7e�E�!����SH9�1��N�sd�A��[���ռ�d񦇱���������n�15�W�y����P"@%��	8v�*��FQ5��G3i|��qWp���T�Ő,&mn7-�8��� ��?�E�k5TG���#올|�>�̸ڇE�փ�n䌸*,���T�9�m�i"��J���;5k��g	6BIW�_6]Պ�m&Z����)�~AGɴ�I�]���X|Obh��F}�D6A��ΐ�p�GW��Fr[���\y���K����-<��<ޚ�1�=�w9l��H����A��
�^t9g� ���D?gJ�d>���Gp!&�eFj4s!GJ�7*w<�R��R$�E��r�~�|���`��r)�vda0�YxlZ ���3��W`�uGrܑ^cbڂϢh�4@��:��=y����6<��7'm0EK�eM���^ǀg#��Պ��.،�z�T&"�m9�u5d(�t�G)l��D=�-3׾�Q�+���,���%%�s���8+�}���7���m��߀�n��t���x��fm̈�t>���oTY��k1l0�2"<&"D�!#i_�2�wGȺf����"�h�8i��S(���������������{�ڼ�� ��X�7ϸ��?��q���~�옛%�#c����&�<'��TR��5�j�0��v�۴�E� U*ŋ�q�f_y�S�|b����Y�Ϯ - �v�t9�o����2����b���}���j�B =ta��� ���}d�}�y�L����2A��t��zy��T���ӣ߰�&�����9���W(�.���=�Ԓ�����h͇`�/�#с��ʀqX�����j��"6���<m������ε�`,��#�6a�0�)�����CY��Z�t}Fea":E��ގ}��c`��(��+!�\�˽<e0���RK�-��Q����[��ņ�T�#4H��*��qJ.�O�{ڥK �d):����,/�u\t쑝��_�M���ev�����(�)���]�,�
+zE[���N�e�b�0���G�^��%�Pg��F<�-e�i�G�1�'S;�0 �4��"�i m��@������r��l�����OB��Wfv��H(V��L�xw�D�D���A���z���;M��oq�sbcC���+:�Jd���)ZQ��蠍r>(MM�i�8�>L�s�84�$�&d�k(s����1_g{]W`�J�MY8�`��	S��ǔ����qO�+RBxo��\�em9Trz#?cq����?i�뉻yY��|�'I̢�$�&��N�Pj;�*�ee�e��>j��$a8a��S���$��P���pX�� ���j$�淹�:��L������D��\�Vi���*�w�Tc��R[�[��AM*KW^��!�@���0R6m��*���5��X�B�q:�!j1{��e�������Yp�qZ��'��x��������?�&�>���-�.JF�Z�߉�NHG��^�UW�\�jH���;�X](��MaqcW�P�H��>o�p�"'9�.|ݬ�v�i8�Q:I��u�[Cm���FKR]O�p��eq���[�`P^Ē��CBPK�W�̲RɅ����G�ϡ�$�ޔx�G3�M�o<;D<~���P��Y�nF�r���B!������d���x�0o�?���&�c#����_4�x��ӊ.Vwŀ��e�B�UK
ⶋW'ys���j~����f$�Z���������3oH��o�Q��]����t���	�?M"�骄:��)}�"��
;�����X%��9�Ҭ��iia��ݬ���Rg{�þ�N����������R4���L�f�>�S;��>X�[���YU��iB�M��Ke����7�6DCV
F7�.��lK?F]j�[_����G�)��R��Gk8���v��s Õ"���H�Z�.SL��Ko�W�o˘Α3]�f�X@ ��b*?LF�{^�2�[�<�+������3F�6s�Qǔ(�����"�M�S%��s��P�mr��}��1%m�����Ix�\W���p���d���vktS��'~#te��6>���O\�T��DM���.[q
����4���-v��z$S�(��[��ⅺkփ_��'[���4�+e�?o@�!��Y�����ɶ$���ez0�]/��Ym� ���^��ix�3. pv�~m�!��~�t��'���]L���p;{EH頚f^�E{^.�~�Y����1�=g��)8�ɏ��2W�����N�������h�b�K!`�m��e��r�y�07����%ǧ펙���9���m�y����`[°�uw� 7Q�+��B�e4�o�$Q���f)4*�F�熂Pt�ʐ"o�F��]���Zԧd���,R�����1"X����AJRS�Hl(~�����G>|&�d��73��u���'
`�E�D��
��"DC�S���tܪ���.w<܏���1��#64���h��� U�)8���b[�i�|�i�Ӌ�̻��^��P����H�;W۳�K�*&	�`3�U� j���J�EV�o�c��ڿ��]A�
�i����U{��c��[�R�o��6`������^�1��u��3^3���	<����v��4I� GV�[��sH3y�H2�t$���J>_CT
@MM��k�{ul����x�1��WX� �,כ�M�,V�U���t$��n	���p��h�O�-x��
�P������S�!��疘;���KΑ�56����H<_�W��2Sz����J�_�K����"r�Z8o��z=WyD�����*�u��*�4�k1��{H$PL�5���/Ǉq�[22�X#$;�s��,f^��0y;K��g_}±����l�g~���x.;���?�����,��cvS�� my+Tz��f��o�6 ��Z����i�=�6lR� ,������t�w/��/24D@*�w͠�a{n��.��S�����p"�i��^��HU?�����`��F��Lj�B'�-��wZ��i��/2Jx:n^b|�b�= ����Pƶ$W�QN�Zq�	@˫J�Z%��j��<*m����0'�%s�fZ�a��O�>2ph(�@���g	����<^�BtXLP[�j��k��f6�Y̮Q�����G�=9G�	D�Ν6�k����aF*9V/��i�q;���'"���LXy�xg"D^T���eF�4�����Z^4 L�N�����*��l�E�ن�,�b/����<�l`��X��.PK�\˲�2�>��PJ�;��9G�]��)��BY��RQQ��3��9�خh\qbe`�j��'��>O#����o�����f���WS��&oI��eTe�F�b�Bzy����+��h����IQSU&/�	C{{����4b+莑W?�$�r��sժ�����"[�O?�gSxb��9�|�d�����F"����`Ʀ����$6{���Kw[�{��y�OZU������V6�W��X�FK"�����&�7R	(r俓�z�/K�krqX`'r��H�����?g[c��=^w�K8��c��	�x����E��j�f��WK�ؘ��I�{*�P�|�4i��E:�Tң�Ce0�ӿJ�27�� �'�D]�i{x7��הi6�Et����%-���Q:�(r��������t��y	d�6�2�΃���д-�4PjgB��C͌I��7�<��
�vw�;�K~qL��J9Z��\,�a��v=��%۶�x?�%J-��thmT�����&*w�L���i�H�\�C���[�0�0`Ry����U������ߞ���u�1�]�7�8X��.[�"��{5�di��,��O�pW�Hv�l�5��U�����3yF�'71A��|(b<\Ά��}W�{L~�i��˾�+<��V� �䯠궉t��AQ���8���\pyd�G��r��/�.�?�9�2�!�/pHg��4�6�'5�;�W�~���R�rl`.��^�ǩiKr��9��H���:��ory�9��"/2����-1h¡���0�\�k+��T�t�E���jq7>�:r���Q=���ɯ��-���"�2�4���u[5�>�"mZ����|:����K7��<x&�EW ���p	�C|��(�Y����N-Yi�>�o
���J�]�*�G���6���q�q#=
�Є�0uX�*i8l�*�Ȥ�l�ޕ��Sb��Kr�P6���f
ݿ�_�{oߗ`�<s�/�p�Oؗ��f-c�f'���l&���Q{�_8H��/��/�hVr�9�>P�m�m'q������_�Jݪx���n���峃�5P]%�R
����)NR��^�dJ���}��U��K�H}��l{�",9v��#�w)@.�Ba���\:�y�^�z۸T�m⮍z-���1Л*�A@Z��'t.人J���K�{���}!�~���7��F�!���O���{�c��hndG�4,]Kq$�S��*�?7c[~}�7_az\��D�B���&��%�(�
��?䀍���r�	�\��\Д9�'l�:�"�ڻ��V�ݤ�Z�1�_J[�+�)�~_�%��(%��e����`�P�f&��+ �����cP�Te?=���