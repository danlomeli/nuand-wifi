��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� rā�SZ )����C.��&0C]�-��[�3�-���+��պݣ�k�J�vo`�A�����f����u�X���v�=�а���]Q�Wۿ�߸�=_Q�X����j>��Zw�K��SvX��ƥ.���#�����Z�0���#7{��\S$��@1I�QX~TQ�E��db����۰� ���>0�%�9�j汈��}��1� ��2���h�G��SeY�a���	'<x�p��k�H`�H�j^y�0�s�78+���ֳ�`�R3dW��_��{p[�?$�s0��#�zS�_��bH
�c�p�IL7]� |����Q�� ��Rr���=��E즕2%�����`�^��l�q-�]�p��jf��Ӽ-f%H���ȳ�>��+���M�71��4_�) 3�46h�rb�J�W� k�h~K0�>P$�_n)���5�r�j��W�J&޴o��$>��6��ŀ�;A~<6P��K�~��f��*I
�Z��}`q���ApC��n���g���3��-�іrO�mF���,�$��@�BI�q�}��Ȥ֐����î�䂧��@������U���vU������ �T#K@f�㯁����|95<@���+�-�)�����K���FI�k���*@�m&���
���ma1[�2�u�I�\�U�yu���o�|��2����;�W�W�}P�K>%5�'�8���׫=����k��,�t�M�0�8]q3���N���GvZ�i�+ C�e
��Ќ�S�v<%���q��e_��
�k�夞��>ZO7E~��5k�TW Aod��eE���G���ɑ-'���?�G$����ќ����8ɸ+ 5ʗ���l�d��,�J�
�^�3b,�����J����#n�zK����z�&��;|�\�^���'e�W�����">�w*	FO�Δ��v���I�h��AF������"�U��� [&y�޿�eox�^�A������Ղs�+<$"�mf��]b����M�m��˫�2��Y��������k)�0H�H���Z�ʢl	�7���@2��'j4i�V+(���9�'<��XMeI fy``�#G� ��0!����b�G�S'����LM��� >���
f�HV�p��@>���VPfD��͍'u�̙��2A�%q}���s���}�F&��i}{��(�p#��ZV�X �@ֹ��{|F�P>�]?t� �Oٕ�ۑB�po�õh��M�1� 	I5=#�$��]5�0x��2[�^���_eL��{�Ҫ����j&#����~I�:*�&��n��L`qe> ��`]Y[�4]���P���~�$�#��0�a"���č.�?>���깠���VD�`l�T�e�m�Y�J�	�wEH��h%��"��y�t������[�w��4*]@��r��mﶈ�zI��b��{�I
h	�d�6ٿ��^�.���d���~�k��`��^� ���m�X�0�����9�x�JqcD�J�4�T�%���#sA��*�@�kp�Δ3��-��>�
9��az١�_BX$�h�0L}g���>�hy��~*Ff�S�ͱ.����fF`6$�U��.�ziImO�C=|f���]�yo!�R� �*���DE��pG\Zx��jP�!$�Z5���Xcy֘t����9��f"�d =��]��x�5�F�����Y�-"O�M��9y�y2�ٱ6�b�@2�I��O[y5O�a�gA������g����6@h:W���h/�d��2��q悯qZS�8\͢K��3���'���	fc��!���!�`s�s��׀���S�,7(���5g�u�`����8hkP"=��d'd����W���@��g���כu�y�c��Ckk{l䳟L����ȝX��yY��&Vd�v�=L�
_�����j� xl-��K��r��ۖa�5�쩌'
�K)s�2�g��:5x���
A���;��c㊾,�ݑ�����u&>ڌ�D|���jP��-�n��3V ��P��B;���:i��4��鵦��M���Zp�����|�ӯ-�����}���R<��*���_��+s���1r����g)�_ӵ�Y�����a=^9hs� �B@j���N�ʡO��7�e:��!ܕ�K����vpn*Ff�L)(�nZxOh&�qM*	�+)�S���G�.������#��-Y�+��C}� �4�pez�Z--�������rP�|*�����O�R��b��<PD�[vB�$��.+��U���t5p~|�ǟ�$|��D�D-Iz0�[�l���^�����0C�f��ss�m~��$���6�)a?�l�sC��Ci�g'w�x����{���`O�R2�R��[�U�|6�;�ѵQ�	�[���S�4�@����4θ�]�����8�߸+�\!���?`��A�8ra��B��(�,d|\/=�埞8��������0�L�a���,u9�=n�����ָ�T��ϱ��}rtK~��fȾ� �Vʵx������6 ���0��ғ��V
	�Dt����g�x���88�_�� �ʊ��`��%��K��1h�WZ�E%^S��%>{Σ.u�eG��<>�b�:���k�C�M�Leܸ�,'���V3��8��
D:�Ԛ�LZo`��t�rЗ�Lt#�!"�7[x7dv
+��#Ҿ�vu��Fi�I*���E�1q����ny�U���#^XӘ��É������ 4^����\�R�%�hW�&,x��M�a'��|��x���ة��kVOL8��ȱK�������η��G�r;g��@y��s���P�q�v�.;zM�Ĝt����EE���Ξ�)�����8m���4\����F�Ɓ"Q�"�΢�uC�G��j$��j���0c�ð^�X=+)9�$���Il�m7��ϖx����U�R�F���+dz����]�c$-�mB-/�	��UeXS��L�h	0����M�<�6x��� ��]�`�/W����w�7j�<J��Dx���dF�KS6��O_����F/�bqr�=� J�0�0�1ow¨,�`_"S�XS�jp����9���u��
@���P�D�i�JyL^��o����n�^�z:��l̯��>6Yꍐ���-x��n%(�x��@�&���eD���93�JNW�fG�4��6Nk��oo�%BKn�c��>5K�5�%�9���_@r��DV猴���g��{Ҿ�T����$�X� Oa+z#��'B�='�k2�Q����r!�l�0�n$^G�eʂnܡ�*.�-$�.���z�A*h�/Z똼�Ǩ  ������-DBwcGk>L���1\cWp�v�X�F�<Z"�@)4O��O����g��$�i^|Q�%J_��5�"x��Ncm����:���{_�A�]�y�L����>��jW�5��AcyDA{������3õ0i���$�PP`_c_�!ڣ��O�CUT���YR�}�����h:8	��ѽG_���Ǳ7� �F^ݽ���n�Hb�h.��?"Dɬ�Uq����H�������&�-���q��7�x%���{�ۜa�@g`}Wǧ�~��j�c���X���zХ2}I+��q��f���D��*��}SR�4*��?��Qv�w��������|�yhf�"b�"�6�:N�9�����w=&=�ł%��i2��/�s�+�Rp� ��ֳ۽0�-^��t�����-�7�BՊ�{\loE=�C������2���M���!�_-��b���}���+��2P 5�H��F�,P\��l���"�~P[+Q����Ѐ�]+�t5�wQ��cx�u�@��I��ώ��m�~��ؙܖQT��.��CtҲ�OR��	C���p׬[c�r�.�M�qf��3�>����e��ٴ5֑�VkI��<;�?(�r/p�;Tfʽb���<Q��h��Ŋ����,�zk$�"���窢�2d!�}���ntc��U�C�#8!p�%����^�r���T]�M8/�A\���.B�V��-CV1D;E��j���;����^�q.C�2�d0Z6���c��E���x�k�%�ő¹X��R��b�F� 6��&� }�f��~�Ƥ���Z�vcg%�~d�$�f��I�L0\�󲓴ЍUpP�	��l���"�ԑ�)[���f13t2�1���ݹ-=���u��#l]�5&�f����z�d,�cl�����O��8N� �W��<��� ������Nw\y��#��<A&�{�