// viterbi_decoder.v

// Generated using ACDS version 22.1 922

`timescale 1 ps / 1 ps
module viterbi_decoder (
		input  wire        clk,            // clk.clk
		input  wire        sink_val,       //  in.valid
		output wire        sink_rdy,       //    .ready
		input  wire [1:0]  eras_sym,       //    .eras_sym
		input  wire [15:0] rr,             //    .rr
		output wire        source_val,     // out.valid
		input  wire        source_rdy,     //    .ready
		output wire [7:0]  normalizations, //    .normalizations
		output wire        decbit,         //    .decbit
		input  wire        reset           // rst.reset
	);

	viterbi_decoder_viterbi_ii_0 #(
		.viterbi_type          ("Parallel"),
		.parallel_optimization ("Continuous"),
		.n                     ("2"),
		.ncodes                (1),
		.L                     ("7"),
		.dec_mode              ("V"),
		.ga                    ("91"),
		.gb                    ("121"),
		.gc                    ("0"),
		.gd                    ("0"),
		.ge                    ("0"),
		.gf                    ("0"),
		.gg                    ("0"),
		.acs_units             (1),
		.v                     (42),
		.softbits              (8),
		.rr_size               (16),
		.n_max                 (2),
		.log2_n_max            (1),
		.bmgwide               (13),
		.numerr_size           (8),
		.constraint_length_m_1 (6),
		.vlog_wide             (6),
		.sel_code_size         (1),
		.ber                   ("unused"),
		.node_sync             ("unused"),
		.best_state_finder     ("unused"),
		.use_altera_syncram    (0)
	) viterbi_ii_0 (
		.clk             (clk),               // clk.clk
		.reset           (reset),             // rst.reset
		.sink_val        (sink_val),          //  in.valid
		.sink_rdy        (sink_rdy),          //    .ready
		.eras_sym        (eras_sym),          //    .eras_sym
		.rr              (rr),                //    .rr
		.source_val      (source_val),        // out.valid
		.source_rdy      (source_rdy),        //    .ready
		.normalizations  (normalizations),    //    .normalizations
		.decbit          (decbit),            //    .decbit
		.sink_sop        (1'b0),              // (terminated)
		.sink_eop        (1'b0),              // (terminated)
		.ber_clear       (1'b0),              // (terminated)
		.tb_type         (1'b0),              // (terminated)
		.bm_init_state   (6'b000000),         // (terminated)
		.bm_init_value   (13'b0000000000000), // (terminated)
		.source_sop      (),                  // (terminated)
		.source_eop      (),                  // (terminated)
		.numerr          (),                  // (terminated)
		.state_node_sync (1'b0),              // (terminated)
		.sel_code        (1'b0),              // (terminated)
		.tb_length       (6'b000000),         // (terminated)
		.tr_init_state   (6'b000000),         // (terminated)
		.bestadd         (),                  // (terminated)
		.bestmet         ()                   // (terminated)
	);

endmodule
