��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$��7�4��L+Q���+2�"H�������v�ao4��	�u��=��d=�>�iV�f��l0�Zs��7���~rM��U�`���e����K%�u��ݒ-� rā�SZ )����C.��&0C]�-��[�3�-���+��պݣ�k�J�vo`�A�����f����u�X���v�=�а���]Q�Wۿ�߸�=_Q�X����j>��Zw�K��SvX��ƥ.���#�����Z�0���#7{��\S$��@1I�QX~TQ�E��db����۰� ���>0�%�9�j汈��}��1� ��2���h�G��SeY�a���	'<x�p��k�H`�H�j^y�0�s�78+���ֳ�`�R3dW��_��{p[�?$�s0��#�zS�_��bH
�c�p�IL7]� |����Q�� ��Rr���=��E즕2%�����`�^��l�q-�]�p��jf��Ӽ-f%H���ȳ�>��+���M�71��4_�) 3�46h�rb�J�W� k�h~K0�>P$�_n)���5�r�j��W�J&޴o��$>��6��ŀ�;A~<6P��K�~��f��*I
�Z��}`q���ApC��n���g���3��-�іrO�mF���,�$��@�BI�q�}��Ȥ֐����î�䂧��@������U���vU������ �T#K@f�㯁����|95<@���+�-�)�����K���FI�k���*@�m&���
���ma1[�2�u�I�\�U�yu���o�|��2����;�W�W�}P�K>%5�'�8���׫=����k��,�t�M�0�8]q3���N���GvZ�i�+ C�e
��Ќ�S�v<%���q��e_��
�k�夞��>ZO7E~��5k�TW Aod��eE���G���ɑ-'���?�G$����ќ����8ɸ+ 5ʗ���l�d��,�J�
�^�3b,�����J����#n�zK����z�&��;|�\�^���'e�W�����">�w*<���=�O�V������0g�R��6��[�̿�r�D`3 (�I����|/ʼ(ӿ�5D�E�)����k�%^��D�	�2I~��|�bxQ�N��.���a����E<����8C�!�f���_ˡ�3
�,c&�Vn4:Xk�7�e�ߏ�5�0��s�l��'�O�24�a�^~]��d�y�לF[x�
�ⲽJ���e�,Y����=ðߢ�7��G�|�l�WEɡʍ��X�E	���&�����>Ԅ�o�Qkd
;��$ڄ��Qq�p��U���9��������� ^�>���Ua���k�h�y�,9m��xHEg��^kJ��3�᫿���$��*�%J�&�D���:�`�+iU������g��J���o�]�7�ݟ+�����3ș$��RO�Bf@��߰
%)G�~X�AC����7�c~Y�+w˿��5�D��q�Sܳ���Y"}翣A�n�.bB�3턪����T6��.i�;�G n�҉��?�N$�krn�{�!Ċ�d�,���њ�Cz�#e�d�l��(���]�8���@7�;���Xz��$fS�mb�upyJ�KY`����B�G�8��Q�H�x�"����CW������2s���N�|��Y;��$ei�p�"�\���V����\8���Ԙ���Y�9�J�0�_t��K�IB�8a�'(P�}��!���*�ҮC˼u��W���ֺ�	��Lt+6��mZ��퇇�L����UbI^�d�'�:5Bu�%�υ�_4�
�k`�^���LN H�'ܲ����������!����V�| �u��+_=wl��h#���_t:`���FۺiMA��M��mHu�}� �6CV�|���+��W�1*�����He�����>��7���Tp[���;������J3z>7��9n��>�4jz���3�0]j�@�>�&�tQ�[{�7����z!�n�}W��y�sM n4�Ga�_q��D���m%��y�Xs�Ơ�Of�ꈒz��hG���R���=:>�G��.�/<+��n ˟b����ܑ��!�Hg2�R�g��\�ev�C�������o�����堵���UdI��w��%�g��|]o��Z�KIp�����OZ��c�uOzYW-٘���S����ү���î&�k4@��=�0%Uس�Bu:��/+�[�f��ti�Q�f�8 �̖��Fd��������Z��G�?��q��(���G�ET\PY�����%�ny�c�H@�Ku3P:��"����5�F 0�U@��(�9n-��%��T�U��o�����%7�u�����p���3�U�ɏ��i�/�4x�}�$�~��Z�#�Љ]��E��p�*�t�S��W ���\�b���9b��0Jw�"L#F���� �Qp�h�5H�96aS*c�{��>Q_�Ȭ!�v��x$%a\�p��J���t�:'��M�",@޼��MɌA����:.����ߏ�P�>\f+�rR���unVM��`
jކlˁ�I	�Եl"��,ʈ���2_��=n� �a�5��wE˖'d���d~���"�
����P��y��!����_պE\�KS��攷�.LSUI,�5�J�_�>�;�v�H�u�d��$� ej5H��:e�%F���4��sH^�NQ#���V,{���>K�:��$�F휨�Q�:�	�S�H�����~,�̖@X�c~`d�/�$gӅt��j�����C���dE�HDQ;lM�sb�~���7��
KC�*O`U�?��B�"ʿ�\Y�~\P��n���E.%��,���l�ȥ�j��A�z),�	E�\3o�y�:���'���v�t�Z����s/���O^�c�\*��!�J"�����!% ���+�Jޟ�hAMEԏ�Ks�M�Dq�����Im���` �:9�Q*�=�кJA��*�m�0b���kPӔ���1ror�Vp8��]*<����e�!���y(EI����N:��R�W�YI��]�Pv�>����۩s�������+�O��w �ڊ�*�ACHW���X�_S/"Oqdc)�3��=�@����\%I���s_j(	X�D����e)~��0vCH�	'b�Q
�>�I��$9�ԋ�Gʀ���;Va��%�{!��t?M`� F���c<� �@f�y�-�yd:�X�[a�(#�	�%��3b*�k�3�����^�4mn�&�^t^`Z{�[�8�����A�Yq��ޓ���ՓG9��w��v^�48�	�^�<!��T�CU=�G�����_ e
�Q��y��ؕ<5�mO�ң�ns@HWO���鯨 3����c��p���|&�9�>l�6�w�QJ��_��.0�#vi�s[r��� �?� ����Ď�����u�4W��C����%�Q�E��k�p�S���}���%y���7��\��*5�ҝ�Գ�:Rӫ�o?�̘���%6\<�ZpxN튗���c�Qy)���s_^K�,(�aA��A2��ADL�q��n��!�ᯫ�o��,{��T~C�q����Z�j�������j�Rt��?�l2���bm���nqH�洏�uG ���a�Ij]�p���Fc����I��ҁ&��~�{��E�*ֻȱ%���_oz�s�55��]3N2��)~�13N�]Pa��`O�Qv��E��d��
��@�j�����፜�T��T�'z��Jܭ���6���3BZu ��Xr��`}�og��-�:��g��L[��^�
 j��&��L�4l~2H��lp�B�t�Ŷ�\�.��[:���6�Jfk��ު뎂��W������U�����(ޒ���y���תJ��M�3
G���>�L�X�l�S	98oV�)��)�U�=(��u�����ѧ�h��|�%�M����ۍ��u��;�	a�\	��xv���=�T�(��]����W�Ex��"�a���)�}�ί���L3���?b	H��a�KW	�RSg���c];*n
�~�X�H���.%Ф\Z+��;�nH����9���\�D�(Ӵ�ۋ�������F�ܲ�"'s��>b�1��~�:r��.*P��Q��w=6%�b�F�g�݈��UU�g��qPr����H�4Uh����M�����B�B���a��*�).)��
g\a���3�I��m��������}��X��#�c��}ɪY�,k��>8�𢶷�`}��k9�]��]�,�ּQ΅��.Z�����3�+�~px�]�́�ڤ� Q�.m멚y�p�@��an�<m�װ�@e%�mׁ4Ҙk�G\�6}e���N���:�y�#���.CS�t�����=�S��\%'�]hMH�E��*��e{���&���~3a����q��=+g%�?�ٓq*�B�S�sƌr�Y�Zz͵nn��_���.��Ѽ��+T4�q"���7� ��ƬN�c����Ou�6��I���a#���΃i67u�����[�hWC�-�m��=����?�pJ܀�>B�G];��/�n��?�B���r��+��e����GO^M�1&�t��e�
��6���f��ѕэ��=+���"�CZ}X��<kn%�Ϊm��:t�LZ�p�[V���]�N��ڰ��'��{�N���*>^�C�*6o�5���o^�#�I\LiCq�#���i�$�Nc��=+a�B�L��2t���,Nn�F��E	�`, �-�����>/r۲��c�}QY��SφA�~���q�?QD��Ŕ���]�W�+�e�ad�� ?Sa�T+���QC�Y�E���_N������$<�$�Z�/�Q��P������_��]^�p'�0�K�zm�9H�RZ
%����0b��� ���ꔶ���!}�p4����1��h� ě�1�}*z�5���̣� ]�R����DK.�	������ƼK��eN	G�ŹiC��	�=3G
S��
p�������6o޷N�C�3���r<�T;��0!	��
���D���0WHK����B�c��/��b˟�0���*>���r\d�B���9c���(�����q6�q'5����Mvߤ{����W�&�?p�	x�%���m�4m		��g�X��ؠ��>f���/n.2t��������.b���������W~��I������x�C��q^���K�4�7:�B�NC�H����ñ7;�[�~���'tӀ+��0�}���������S�aP4S�u�D ���,�Fn�V���҅x�y�"�U ����6�QH*7�^g������?�<�	y�2.�;���F���T��!��z�[O���4����Y!�} 1��(HD:l����->���+��8mLc��*��3 �b����8��ow��cZ�����ӣ��v��v� ɨ7­�5��a�&*џ�H�}�`L�7ė�ڵ�Yy�H���Bw]����\�֎j)xb#�jJ��#��E���R�B�{��m�hΦx@v�!���>PW�ν��Q0�b;;�C�M&�-Ņ�����lP-2�9�VR�������|���^���R����7�o��bu��h�%U��e���3��瘞�Gz.)�+Y~�H0�q�Ʉ���G���a���F������~`V	��I7��8�Lue.Lx�,��(b� ��D�D��������Ρ���t~vj��/R�gh�Ԡb�9=r�m3��H����[�s��լ��߹���X 	���+���7a�p�yOƸ��Kf)J�Obv�s�Ҡ�~F���v *v��&m�1mqz��f�~ҫ���k����i
c�Su82��J9�%�)���oO=w@Um8���f��@*���v��?�	d� ���C��9#ߚ&m��$F@��kd�t{�jn\��E�&�@^ʄ�y�z�C)O�%����a
�����<�dr���7�	��6n�7X�&)����k��<��8�
F�ͽ˟��)�2�'Q� w� ����JYm��͓�ns8�g(<�gN�e ��b��N�p����IHͥr�C��n���J�����ŀ��F�e�/�]0��, uB�rV�����<2s�.DdՁ�J�����b����c���e�P��]�n{�(v:l\1��>�w�@0�C��=���5K��s܇\UR��f��I��G�K��_�����,�`&����<���
�F=�5fb��zځ٥��d�V��o�������|�@�b-R�_�c��=�!zpx��:��mu+�+ANIt{	�#w9~��zZd�G�U���C�߯&�?��9C=_�^�a��߇0�l�EaB�u����R����(��<j;-G-N>��Ľ8a~�M\�:E;��Έ�0Gc�v�jO/���Ί-�B���8��� �a��]ˬt��$hU�r�L�p���2���m���x9��G���&�\�Ⱦ���R�=���/�bJ! �/�5ń�]��C��͙+1�FѪO��=���P�@V/!�p�֭�v0n�����o>foʙ��2(=�&���	4���w���jN�ٝ'��#�ymuM7�7�<�h��� 'WV/���(6����/�4K�͍����P*��v�����M�_�z=�|?v�7�T�&�ȅ���NN������'�!)��%_2�C�hk56��M�}/�ע0^���FT�Z�(��u������$�R`wܬ'r�[,B�6���Py�.\���pDo�"��7tǙ�j8I��o��u�.ƽ������8n�� �	O*<��#���ᆞŐt˚��|�֯�,$���%�g���8�+��Pu��ۀ�r���u�o�Pq�Ϧ�-�|J��߇b�'l�W�������C�`�ؿ����6�$1׀/������!L��x�k�ۡMMM�<��E�~��SBʐ~?��y"���n֭�/٬"%g��y��z1^�[�53�s%���b��B͈ɣG�ٙ����T�	��q�gΠ���5����߰�xq���O���-
�P��|�R�T�$�?�'�/Y��b/�>h��lz�:o�Y��"�b&n��WO��N��?nvj}��`o�#���q�R:!I��B�t����?<&mW
��(��id��h�6)X*��>�2����hl��:K	������~�J�72i�KWϥ��C��1H�~�n'���+�����~YL=o��b���!ڏ�_�qm�x�s�z��9blN�{O�N������v�>!�ip�<Jȑ�&v�<�D�,Vw����-᷿����/���֧�@�(�S<tR{�:[���|-/�_�ʩ��Y���ae.V٣=�J�*�!�<��������n5ȑn]�~������'JT���*�I=��v���e�~�*���ø�[���/��P�
-��T(R�δ�E��{'��u2�ʻW��u�%o҄y�n�P�:�!΄���\���2�j�&�l��g�7��� ���'�N�*Q�i@3x����Y��h�؈��~9'o%+�}e���J1U�G.�[����6Jb�G[Y����
�P��僂���?u�{��dB�tl:9��4��E�4£��9�^�sS#�wՆ���M��JLv�kR_57�ܤ����!��xE�z�M�o����t�eWk,�������OA=�y��5ODi��m>��?�g!�WJ6�n��~�B�����Sԥ	��Z��t��_�zf���/��(�=}�ك�cY�r\;#�u��u�����<"��o�n���?y���X���A�͑`�)�Y�����H�ܙ�(����'\"sd�4@w<+'�[p�W����K5��R�!{C b�{�5���&M��䵆�}��܉�'�j��ˬ(��^p8֜�m���qJ�a���X�{cbN�o=�n�i����ۜ�uڤ��7��f�:N��xَ��R��6bm�Ho�.6��[��� �_�y��s�Gg�T��u����x��!�Q�0P�9U�,�YU��������k��R.��Y$�Z��R�y�G}���Gܴm؝��Z�e��S��&0;b`�ɟW9ˠ��(�! :s�ė�y��"ۢ"}z( �(@��f@t/
�hM\���H�X�Y��H^��U��������=1j@�l3&��I��V�b3�v����2(
���6���{�?�]M�u�b"I?��8a��¸L~��%�Zorร��-���k_E�#�I"O�h�4��b}rx���K1��Ҿ;��b�L.��H=�3m�&�-�C��b	�|>7�Z[��t�C��e!E��c?�?�r�2��B�OE�	������sc�LÑ���K��#k�f�EG������b��$�,@,y���'iv�u}3�`��hT\���jx�M+!�j$�����P%�S�W�m�c������BACh�i��IA�9��#�6,�_2��t�y���I-z��lF'w7]0ʀArH�׾�pι)9��``��vg%`��tk_n.�d���H�S�Ԥy4��s�����!�crT�3f�Q���t	��T4�{�1�M�G?4�lQ�b���t�aw	>�?)z��e���;%T��S���wZ
>( f�w<��1�,y&��M.�L�Yu�Z�J���|H*�������h�Ӳ?=P�-�(~P�E���J��vkS�yR�y� ��,�9M|Tڊc��s������c�β#�`�3�.�-q]@��	���.�-2� ���������G6Y�*��*	dXx�}J��$�
�.S�V	�*��F(�bIW�ht��]۹ܵL�@�JuL��7��������C��;�j�.����O:{^dUk�Oa�(��8_�0k�Hp��*��6[�Ql�j;�l�L��u�<��l�ec����v�2��3R�ʔ���ǽE�3᭽��q�kJ�p4\t����ԟ��6En��xsQH$��~ܸ��� ���� 2�{�r刁��m�c@+!)k��P�k����N\BX<Ŀ�Q!���?!�t{.~.�Ik���@B�C*��|��S�~[�_�:{�:����L�5F^�*-q�$�7�kT�t--�<��	��CV�7�Au73�T}���)��4þ��X^:@���RF���J�����P:�F����5G�c�pR���)�q�B�a�N��f�iA������
%��R�OeX���Y���`a����YcM��桕��%�����?��9�0an�)�(�����Äک�e�?�Gm���#~����dc������ +�e�hU�#�D��Շ`(k�+��90�)���-)զ�-��r=����� �A�����ؐ?�L��!V.�<RC,� �#��q]\��2�ςsiat�g���^~djt��2�s3�;1<ʩ�Z>�
�M�_2cr���@���P �҈�#�ҔN�q��=<�4��\���?<��Q#��*`�z�q+��)�bX��L�)��^3GQjaELA�X@
r ~��vR�%���#�p-z��§��������z!�[y��PJI����f�S���2�$.��qp�������	U�(L�_
�9�k�2nﱀ��W2�,�ez�0i5��g�0)q���@�˨���Zv멦b@�7E����456�;�"ğG������u���1�� T&�<x�24���Rm� �WA6��e�#��Sa8��T��'��A�[8�NT���Jr�G_�yHL�җ|��IUi{����瘻~�c��d=��I3��ڡ�Ǟǝ����À"�r�GPQ��ǟ�a��ܠO�OD�6��Bu���6��ϰ�5e��k��E�j+��(�e�<+%�P}�qY\�+n���K�2��:����EH[�r���d=ʃ��_j�b.$�v����z2j3�0�� 9]J@�w�#j����5�n���rz��$�t��=3�[��3:�J1�I�~�>A$��ض$^\�$�".J�}'���X��n�{/����fN���*��Ӹ�R��Ю����H@�
�s�lx9�O;X싄�q�%0Q�v�*������]ˡ`Ej�0��&�ue��_��hp>�sU�Я�Lc&x47�I� J��	Ţ��_��&g~�X'�����c";& �(g�����ebUoU���s��4J�1�hw-�e�˔�j:������Sk�Z��`�Ώ�c�g��aϮ���cʏpꉦ�&�������wy?�T��u�M���;��E{����N��C���e�M�z?[��cV�!1�c�c����L�^�����>J�����k�[�|�e�f����[�����l���tH8�Z������Q��T�^^�j}��9{~i�{��'���_L�!�B`���f,�*(��~�qPKkV7�T��1��9O�������`��Rŉ2q���@	��Չ@*��9]ּ�V�,`|q����ϧwzS���+������g��e�UmU#�An�դT�k2���Mz�8΅Q�P�L��qB7p�a�¦�ޝR`}J���^�-'����y�����1�@��<.������B��Ԇ�ER �>۔wf���P����
�"gA� C�q��'��s�3r�� ��f�Ě�
bt�!���7��܄���y1T�V�oU����%%���T/.3��'wzR��y����{w�r���I��*�+�"""܈VN2�����G+~%�^���a�(QHށ>�&��ٱ����yNՊ��u�d��~>~�̑m��4�iuR�;w���!����I��'^��I�
+�N��E\O�0h�k��,�Ȕjs���F\y�1���ae�&�#�H�:ÿ.��|<S8��cS��YL(i��O��S��w4���!�;��#7��Ng��]�N1h��Z�<��������A�����L��F7���U
���uFm-l˽4�ȭg��&��("ӫB`}�H,�"����	dJ� ��2�$ꬡ�46�o���^4I�y��A��l��ŏP��A��b�*��&ʂ��K!���|⁜ ��S�"~�C}����R]�>@˵(#��hW��(�҇t�ı�|ߊ�HR6��#�ˣ0�~ޫ���l��O�f���U�������D����p�Ȟ��y�J��g�B0����O�7�׬�]k,����G���ܰb�y���Z��]����b4��4O���Ge{�"�A��e3ďc̕��k��1YD�A��]�k����sO4?Օ,��&\ݝ�~6n~R;�k�]��K�)�������&�P����/��刌���c;��?^W/>иIX�Fc_=���*bO�����1l����9:xN�����������ʯ����I�\�3N%�0N�aI`]o#Q�^֊o������B���|aG�@��8LA�p�fx�'�u���Ch׬GI�69l$ROʎ;��V'�����<Q�s��V�f�x��~�V|l�:��KP>	����4���%G������F�\�n�[J���ţ�<Y�A{t9)�����8��~.ģ����I�"�w�j6j�����W�}<�+�Y�N;
H�3�RS��=q�R�r�W��{�Q@.E7�.�'�0R��66��Q9G��O7��xx�[ɡ_nZ�������o�(�痃��m�����޻8j�e�W�����$�6�2Үa�����U/�`"�C��b+�E��O�b-�۳�(���y�{e�𒒴��X�����/�nTt�d�ľK�����2Cى����q�`9ӑ����S�J���H��s~�L��D�s����ѭ{���B@�������F.S��P�i�+����h���@�6�����)����g��G1��F㘫����$Qi�1���"ԇ%����G&��U�x#�Q�4H���EO⡾�ZA��`��K�Xe�A�VLG��E�*�qǝ''go�
/��wӀ�~뢽*"�J@{�+��}1���.��Dw��A��W�(/';I���U@����׸��x��M	��"2&�3�� n�Ίց��$��
SP�=S
?�O��6{U��dN�!�8�;�̰��J/�	6V�pOE)�E@���'����Kgv�O/�Hњ�߻�?b�����5���Zi� P��C?/�!��|��q��4R��X�?+��p�,�C5�c:{�!Ȃ�L�F줭�L΀͏=�����@�0�/�ItGy��>�a7}�Գ�=�9e'�k�R\�(&��:H����P��b�g��G1�僗ݶe;ު7��4\X����F���Q�:��Vz���N>��U��Z������������<�IS��q�-�2��}���:����t�V���Ssi���yF�9���]�㞰�ΎW.ԤL�%{Ȕ����AHV:��sNn!/�n\\��u&A[ݧ!��ϑ���7�=0��Y:�9�z��-���g=�O�VZ?��qG��'�b��Q�� ���ZO�/�%g���0�I7ʑ���u'��J���@�f0�]sը�S�	D�XV�ׇ���U�>O�Z�`�e��d�Se�s���#[�NY���+)#�đV�謗K����&�J5>��6�ז��8<i�=:ʸe��}���3#������gE��}o�vg���w�>Z_WA�ϼ;J��PV.w�!>�w���X�}4I1�
KEsjJ���8�����wk��B�ue�g?���C(���.X� G�-1wm��_�I�߹JVB�.��	�F��?(5q��g�ɷZWq���A`���]{!��i�&91Β��:*4E��/m��|�W���I��G����,ۯd���>7bB�r�b6���2E�8u��u�J,����{����U�jQ��U��
�ܡLg+�W��Mk%J��ո��@�4G���3/�>J	:��"6����>�6���<������d8Ċ�cJ�]�I|��[�Zl�5�W��e�Fx�]��<1��l(:nAe�#sޭP�n�7���L�) �cfF��Zy���S�n�a[B�w+t���H�6xp�@�P��'��-V���9H�	'�#��O��dL������j8F]�կjLBd����F���,��?���LBu��f)0�~RހHFsN��3�� �d-�0�u_QB��}~�L%����۽��C2rd�i�@�F4�����7�����I3Co�]�^C��^�1������N�����xy��q3N���XinG<�~�v��w�]�����l�	�,�QG�����4|8��EI���6؏�4!6mEIO�isu�
��2 ��l|���f�KoQN�i���.��?�.���|1WF�"2�u�Y�a/8�	�p<�ER�/�"�@�Z��!�s�A�\CG��5�,z�~]����p��j�@?�)�I�C�|�y��ʇc�L�A�S���3�-��S����f��{�]O�#�3]]��D������<n��x`f�x4������=��υ�Ȕ�f�X�;����.�"h��;A%�9���cM��������49�|x̘�_���
G�2��~�����S�۠���n�;a!	&
�����wP�eKJ�,�"YeL����$X�.���K)��Q�E����� Av�Eo�{�ɷpz�}������v���f�M��/����&z�������!�!P���&��)zŤTZ$�������9K��JP���ݸ(���W#����������1��Plj� ������++ʕ����8 x�6w�v��x�p-8ͯ�wpoK������:�S���a�-���Be�YO�� ���K��=3V<AQ)�;o���|^V�U�%":с �L��#��껂Y����n���ܼz+9	i�<�}���p�m�V��:^���)�ۆտ�Y=�dQ,p+M���ܕ��8Htl��/ܩEM��/
W�sX����u����%����ṵ}1`�sz�$�3|s2�I��yL	�(ʳ�B�K'��1��Ƶw�J�u�P��E(�	gE��t�-�av���ο4���(�������	z`��~��;z��p�+P�H�w?*A��r��+�f��*3m���=�E'��J�r��Ʈљ5t�pB*D�4�u1�ǳ�t^Y��0�r��P�S�͓�H\�&�d�F��8cy�u�����Tm�LHkN	B�#�����tsol��D|��-5�R������Y�ܚ��0��>@�	-��S�������'Z�
ʰ﫥5<S��x�Fvʼ����;<&Ox�~���nc�b�84��ό�V ���;O�7m��,.��\��:�� v�)b�a-H|���~�@()b�*�����ۦq�3�)���mC��)�|��~)��M+��G򂽓P�Q��(��\Iu�/D����kz�"��D�ᐿp�m�OlP)�D��?]���<0��Ëin^2_�_1��yT:C�7Q�m{f$5WN(�F�|�L-�m���4ː�-�#a�쐩V�]�QK�>5�8gD�%}��#O��
Z}^��:Ї��q�?��&0EU��#�a�n�CH�t�}��� A�;y��A�u�L��!L������U�"Q�3,� _��b�:�؀W�,TAv�RT��,�:�W�P��ш���pR��:n��-�.��
jˡر� m��U�4H+J�%�?-��F�
��������F���W	�?ϯϧm�p�eJ�u�gd��pW ���s3fL)�J뉫��xh��#~��Yz�+լu,e���f�Ƒ�	?/���d����,9D�ʌ
��"v�2x��{�� z����i�kA�;�;p����J4�C��gڐK��N���A��|d�r{��1�Ϩ=#Se�#+���Z��+�WV�G%��ߧ��о@�y>Oz�ȅ
��/&h�[�i�N\�zռ���1r���ݎ��hR�R��������#�� ����vх^�a��^6�K���u��9ɜ�;�Ɵy(��%O��Ώ:3ӛ�kk��u�9�Yzg^25�Z�M�q�����n�O&�ܥݚ�?$y�ɇ8E��Ƶw�2'�%�_W��Nm��S[`�fn��@�W��僣�E5Df獕�D�)gi{��Flxx����:�����^��I,�q<j˿��[?9�3\�����o�By�W47�=߉ �x�j�)1V,�r ��	�D� �KRﴬߦn4��{m���"
Ε4�������GB-�yk�����}v�s�<�٥v�^�Y��՘Ipf��2�ͣ-�?�&JUe��5���(�ؑ��hQ�Y_#� ��'t���'0am�w-��{RpTK	�a��L ��Z�ܬm��2���1@<�HchQ�l�-"�߽��M�9-���,�|��>�;H���Q�����8�� �
�\�<�G����%���S�#*�8O|]���ICI� V��1�(�F1&ùL��Eyُ"{{Rhz�o�)�$W��nס~������ܺ��)E=�nC�!c&<��*INH?�xf>�1	4M�l��Z���|(�y�N ���)�� r�H��h�4j�AH=�zY�vk7���N�9�V�]���۸��	6k�ݱ���=,�:Ο��h-i�#�l��+����L�B���H� ��N����v%{�[�q4��l�����yo^�.7׺zMy`� �-V�j����[^.�=L����b�j�!.ooO���o��tK�>v��m�b�y�׬~�?�q��C���o@">}�4��f�M:⼽�F��]����	�.�Jv�!����E9��:��A'R�l���w
B������	�������+CEM�d6����)�q=��������@̎�"�K��� J�S!��/���@�|�ym[�C)��吾�3�2�����j�~��|�����*Ft����r_2����V�
��G�8Z����.ҬTw��=�cQ�^:f���~��v"u;���'����R���Ȋ
�5	UD� �_�� �٬�%/�uB(�	��5�M:����ѫ�\�ݫ"��kiҶD�a�=lŰ��G�#p���� �W�6�+�cB�NN�"����'L3R����*wH���}�䷘�8�f�Z5/j��z�W�5c��]��>�ζ���$GlΌ��!Iyw��������MiK&|��E�42'��-��'�!;Q#���+rH�]몺�N"�d�oC@%՝�w�mB/�kz�ݢ�C.b�?=��.r�No|�vw�=)��`��3����`�2�&�>�5�e����$B��[�g�W����s俜�������Io��%�hǽ�q���5G��;����m�0!~bg�}���=�&Ѡ�)�\��L�9�aJ����0��[�@�%ؐw��fg[b8�ﹻ�',8 �C*A�eڶ-/��I�)�5�J��Ҧ�	�]��2�Bb�4��Π
��'j'�s�"A��Ś�#�l[��0�>&5��@���-��7bNnxx�O�;�P�V<����s���?O:U`�RQf�1Q�_������L�J�K�����q�0poM�R�e��C���w�^e��i��v�Q��z�s;`#��]�P�y��>NB]_Vl�݋�C��h.������L�a�Ny����Z���9Jo��yV4!��*Um6��3��0��X�N
�����4����r�N�R��� 	 o�]�,(�o���R
�"�Α��}���PjVyd��0C4d,1�a.m�R���5ԫ�5E��h���Q��]�;�2Z�`#��?S�q�Jt��K9
i� ��Z���S�.4��
�_�&���#�9�R�)����]�7�e�6zFɐSeP���li�p�of�Uh�鬻�O�^gr����5�:����J�n梯
*������d.[g��b}݊ZT�XTՕq��g ɟ�\Ie}�#�A�L�=	a��,�g:r��T�D�H,+�F�a9�D�vR�"�R�Ǖ��8hJ��eWe,[��2n��]��P#���%��o��MQ��pJ*^�?dC��AЈe� h%�����G
Ơ� �v�7�~>�R�c��`�"��N�Tk'�*���១�5��>��£�9,�h ex����eO�E3`�Ty�>=ܼ\j�W�uF�N�?��QҼS|��JܬF��8��&F��E�P�'� ��c��W)!�n\21U?7/2Sq�Ѿ��u�`+[M���0�8QJ�C)����� 0d����=P	��1�.�K����(�R�1{��I,m5��(�c7���V`�}��}�%6��l��F��;��}{?����*��K]�I������#���1(��B�:��/�KY.*�!e=`���.y ��>��VT6ڸ����K�1�C�`��]��=��T*i��+MX���#Bl��i:���l+P��65������q�M��%�GB��b�Ю&�N�T��vʓD&�%�v�E��Q�τU`�������(	�g���wZM�u�u|<n�g��>w���)�1��3�R^�7��A�az2�ʿ9�1؄���\�<�g���w((���+]��=pЕCxg�ib��;���JfQ������dK$��m�<����0+DϬKbY�=���bV���)�1�⋲�HUK���A��Ԍ�zA�Wmn`��}t+j# :0�9��:��D��^3R�����Xx�0�F ���I�u��g*ɧd��������=�-��yQ�g;u���"X�=��0")�;д��]���4�%G��ҸØ��z�)�
�Ug�g�(�Q�������*@�]3wн�@mORU.4���s`��7�ٌ].�^�Kc�Q)�p�O�YB̋?]��{��� �zfJ�� �=j�!zA,�9�ёp�΃��"��6?�|�@��QD��2!�:����cc�K� �2Qh��d�GX�`�xHM�f')`<����V)�A�#T�Ԁ�C�x���٪�@��	��8+����A�-�S�3c���>eRbt�����<�����I������ސ��>���c	��@�l:����F9��iv�习�0���w��}���\I��Q���*c����{%�T���t��l�uWN��sl��:�2�����0� pd�qgyk=�Bh���_4�O�oT�e���"Io#Z���?��2�����Z��z8�k��t��f�O�@%v�ĥQ�cTV��(R.�Le�����q�e��(��H�����#�#���&oR��9�+�SA��}���tN�G]�H����){����Ao��Y�Ǒ�O����Y�&�O��;���V@� ��y]�?Dr�����4Ӌ�/�B�	4gZ��X�BI�^�C�3/"l�uݳP�	�������U���DŔM���`��SbB��QZ)n��E3���.��uk��&���]���(������D�'{m��T���I�6Bj���A�5��b�+w�FYQ�&$C�t��M�;�fry���d�e���@vu!��������"���5�2����X�H5���d��>�O�"4�/�Ql�ڬN9k�l���){NP?�t��۵Xk3�1:��N��<F���1���Y4Ӱ\D�~6�����4$ ,¶k�P�h���%��Ga-L� W��ѷ��xi[��)^��
��Q��H5��r'_%̈F�G���V �-j��M�'߹�'����7�fm(���C)��+I-�K���l_���#:�N�����cc.o��I�����_
���^mY�w��3�m���í���~0"�62Ј�h�!�-�*c��mu	����1I"��#����o˟�s�)4�l����y�f���������>��<�b�lxV�.�=�7z8p��7��*��yICn:ŏ�I���[_��f��b�>�g?��y�^W�L٘'�����=I��,��'�'�4y3�s�;�۸����V߰�`'p��Mk�|���m@Ђ]QI���B�%�_JkܚN750o�����4��(����jN�ٮ���لv�e@Cz��4���8��_A��w���6�@T�<�U�'E��	��>>����'��'c��K�n���`Z�6{BB<�����~?[�j�$�|��eDR��;��"qgd_� ��=M�L-]�1�j�G[w� C�>��_7�t�뫓�J|�?e��^�0��;t@��[+׳��^�� F���^KK�qy��XA)�K��H���rq�|��bL�7+���R��䆶�V����LU��T0U��	����j���bX �kƤ�����oQ/޹���"��G	��r�+��ٞ�GM4��8��$���*3SC!߂���I���w�-g�R� RD�5��,��(���q�-c�c�Fq�"��+�֗�\��ߵu�?'dTX����]��3�����=�v*��E�S�F��EP�?6����Ģr�&9�Z����<Q����N>�
����p̂U�
���$ۍ���ri?խjЄu�b>�~�L<(j��_+r���=J��&4�]�5�3��R>!�>�S��^��6l�����J~�P(.zw77�S뼐Į�F��i���=,���ʺ�P^9Ym��+�]Z�2|^�t�<,��>R�{���l>�B�?�Lثr}���}L�{S�0��5w��׫�>Y�t�b�BV�ֈ�?�����椳`1�|^-aE���'KD�C�b� 
+���}h�a3��f޲y7%�'蜿'��'l#v�t?v�>�;D�؃���o$A����#t_%ŵ��K�+�XJR�n�q��G!�U	�`3�ci�C:y���f@���p2����o|-��ﵦ�}۫���킫pz��a׼�;�rTV�<w�Ѷ�+���e�;�u��Z��4I���Xd	F�����s�l��Y�A�����0{�67Yq�*�9�7[��}�}����R��c�E��y�0��NH���g�aJar�o7�����d뱷|���ѩ'�9��%}��!�k�3>op�,6Y ����"�Z���F�֓�_�� ��1"�DBK@��T�d�B7K�@�W�N}A+��W�Tӱ��=JC��>���	TI<H�DJhF��s�\\���[����yvM��l4�h$�}�P��~�HKK�@W|�C&������pc"ݨj��ha���d9�"�#@ŝ�$���-ߥ�Բ��v��"���0�����.�%�q����2�=	V��:<R�+*�q�6K�h�%�mo/šw�tT�8b�G�����?:Y ��n�䐐�Pۡ1��w�CZ��/��٦i?#�p�/��"'�q��� $e[ n�4���jݬS���il:���A�����-I�������!�@3ܽޏ���#� O4�I\���P�@�-M�^|��v�YU� 28sA��ҾӦF5���FM���}�M%e�G