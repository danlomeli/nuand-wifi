��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� rā�SZ )����C.��&0C]�-��[�3�-���+��պݣ�k�J�vo`�A�����f����u�X���v�=�а���]Q�Wۿ�߸�=_Q�X����j>��Zw�K��SvX��ƥ.���#�����Z�0���#7{��\S$��@1I�QX~TQ�E��db����۰� ���>0�%�9�j汈��}��1� ��2���h�G��SeY�a���	'<x�p��k�H`�H�j^y�0�s�78+���ֳ�`�R3dW��_��{p[�?$�s0��#�zS�_��bH
�c�p�IL7]� |����Q�� ��Rr���=��E즕2%�����`�^��l�q-�]�p��jf��Ӽ-f%H���ȳ�>��+���M�71��4_�) 3�46h�rb�J�W� k�h~K0�>P$�_n)���5�r�j��W�J&޴o��$>��6��ŀ�;A~<6P��K�~��f��*I
�Z��}`q���ApC��n���g���3��-�іrO�mF���,�$��@�BI�q�}��Ȥ֐����î�䂧��@������U���vU������ �T#K@f�㯁����|95<@���+�-�)�����K���FI�k���*@�m&���
���ma1[�2�u�I�\�U�yu���o�|��2����;�W�W�}P�K>%5�'�8���׫=����k��,�t�M�0�8]q3���N���GvZ�i�+ C�e
��Ќ�S�v<%���q��e_��
�k�夞��>ZO7E~��5k�TW Aod��eE���G���ɑ-'���?�G$����ќ����8ɸ+ 5ʗ���l�d��,�J�
�^�3b,�����J����#n�zK����z�&��;|�\�^���'e�W�����">�w*	FO�Δ��v���I�h��AF������c�' �J=)�&�/�K�d��dG�4D!?�����t�"I�Y�ʫa����e�N�llEn���AB����~���#�r"��Ӡ�.���i'�a|��ZV�p��VtF���L��g-a�Y�S�'�I����`;HY)|o�?�+:(��.l-��J�<��x�iQ+l���ޫi�q�g��}��5�y�a�#�g��J]����_+BY���B�OV�kE5���toF������d @���ƚˍ.}UY�lb�V�'����&P�T<u7d�V�ȋ����ԭ![�H�L��´�!���w}ҳ�Z�?��3ǳno�"E'������o~�>���Xz�
-(t�(������L�צh��a����/��PA��m������4�Wmſ�nFR����`wW�mmT���|ű�kmk�뉤a��p9!����^��yO�\G�("t�~[/�P})?���s!��,�O2x9ھ!�-�ء�,���V0G0Э��('���+<���&O0���	D9����D����p�؅(����Ewg{2v��͂���S˒<�����*�$}����Z�L�~�4I�,H���&9v/RG�X�;��xk)��k!�+�&s'��g"�?ɢ��i�/�C"��CbtC_b�����z��'Nv;
,WV[�F�rH�9�P�l
�>؜�]�L�p8"b�\7U��3�[12�a�����b:���͂�ӈ�Ι!��?�_������|8�7��C�Z�sa�����,Ca��.V�y,�������������/�^M��A�c��5&#�1�����E��P~�Z��V3j&�,���S�����ߢ@�fkzgMW;2�#���^�4^����n͚�#EYTu��1'pM�Aa��A��֥��<��Wh�d�T&ʀMp�P�����Ih�&8���N`ӥ�,������?R���Q.��l&�c�"ۂ���x�B�h�����;i'�`V�'�Xb���C�~��3�9(��(��Ẃ��h�~��L��n��ˁ��X]�؟�����fp�o�s�͌`;�[��j�u�?0jR �1O�l��&���n���+>9=[#��ڬ��Lsu
�,ⷊoϞ��B
�� ����-�$�d����6�ꪬ����3�e�+=�O���,<�C�R.�����ߥ��*w'n".-�6��<�!󜏉A������s_'e$�r��v]�t�")�Z�h�#��Ax�+��UG�0�_B�ŋ�Gb��I�5�q	v��H ^�D��4�����C��Y�һ��jg���B1�L��uN8lSy�]�C��>���rd=�����5X� =M	�fa�����b�1)�z0ט�z���w�������$ZZ�f����=u���±����i���o���cju���N�}���r�A���?��4s�+Ƥml���@#�Ǖ����i�+�c��Q0��	��xFT�!�p*���Nj|go���d�<j�����u���_���6��G ͩ���:A��z�z+�y�:��D4Pт0�b�c&jҬ" �F�!�b6ɢ%#,���~���P3��h�������AW��,�K�'�]xV $��S~�����3�;�M?ܹF�u�a9��XFa.uZƔ�ab��&6_x ����L���:p�/c	�v	�ْ����2�~�ۯ�l��2�����;7>�������CL�� ��M�.0�Ӻ^�o�����B�H*���]�Y���To&j�2�8|�H#dY%�AK\��17{��b�~?ʨ�m�(�U�9�a���-A�M���8<_[R'�k�|{����	�^h��G�b&G�X#֟��s�n�ꏀ�)�ql���N	ɿ��Y"��J��pe��"��̖�[�=�P�áj�F��>pHK)����#��Y�I��PH���9L������Sߺ�)��')�a^\���ȋc^�P�G�yY�a�S�Zp�u[V~DYg�N�|���1�_ +��A��3���0E^c���=:��+"�̚�l^�3p(Ӄrc�o�vQQ�PR�ϝ@M�07j��x���x�'�'�Pn�7���>�#��XSC'��Mb�t�Q��E��F�5aw�F�C�Z�ūj���=Yw�`\8�ǎ2�MxC��х&�b�}]Æ@x��j����&IVDQ���<!槼s6;�nk(�TVǉ���H�{���t~�B4r�厬@wW�ȥ�<��8�����dD!K�0T���dʠ���t�'0?,8����y�N߯�ږ�lQM��������S����{@CCd�l�/����,��:�t�
�9{5����� �$�5if(�	-�r%����	���[�2��'#?���:{���F��m֟�-�~�_V��rZ���B��T154\X�]��V��$7q42��3@�� �4##�X���d��\`.�T�z]!}��-tᶱ�t��x��� ����3c�msNqFE�����Y��֛�z���2s����i*�����	f�5��]ʋON�iP�U^�l���^Ȝ���x�ć�O���ȐH��|}u�yT姳vW1�Ӷ>�*ƨ�����OE�A0`Z���EZ����y'W�!����9V��"�q��a9�9/x"R�wcD��M��R����@գo�h>�ﳙ���[���&:�7�ċ�l���.��4A{>���'Y���h�e±�8�����{�~/�#�&jp]�d�\mc:B�m���WV���k�Sa�4e�[d\�o� !}�u��nc�u��9��]�w,n\��c0��_ɛ�Z��~^����n�[�L^�[��]n�ɢE7Hĥ�=ٲ����%�*.��톫���c�5�,ܟ�6�<Hі���f0���FI}��k��� �:�va�|H����'�SI�Ōs�3:53��"�?��%x��t�Z�0e���@�$�Q�3���0f������zm�0���h?	i���z@�1I񯶩Ҡ��*2u<��h=d�o#���b��w �R��SZ��!{�6�T�wP�ȹ��$v�YX\�t
��~��\<����M-G�L! �]ƈYىDW��U��Q�`�Zrv�v%ؒ``��J���u��l����	5��q�~	���dK��������;��d�}�@+G�A�^df��7��(7=~%��t�P�ά
i櫨�NOvK,�(����æ1Gr�+'�Kj��1���4�R�++.�T�kU~o��NŻrp�C�Y!�aJ/nm!c�XfL���j�NlRh��6_���E`J���>{���;���t�,-*�n���
Lj�ȕ���B��7�6|�ٛ(2R)��T�/�D�����_L��AR��y������Q��2B��hfD��9���K-��!A��������{�acLdY��m���?�`��9�PV�G����mS�A�����(F$!�OҕYM�[52���Uͥ��s�
�K���8��`���-ڱ	�;*@���͖,���r���2��(�BT��ϟ_F����n6!&n}�Ȅ��n�a|�}�$n�?ᙖ�eI^�(�.���^_)�JIsj���9��a�|oH}Aon��#A��Q��9�Xh���!�S&���g���f��lN�Ƿ˰~�X(�����w�ӨHP�ZR(��%~Ki~��A ��ߔ��ѕ��
�d	s���IVa�7m�B��Y��N��אQ3s��b���x\���q��!��*9�ϋ�Ft5��_�W S��(�2E�3��L����"4�"��k��)6
��Q�:I����J?�q82*a�v����`��Ma�z��o��}�����&����˲}�B��A�[�?�b���@�;�ϭ�qP���J?�h�m�Nx��w
�Λgŭ/�ʈ�k�L��Đ�=jߗ�����2~?33�h^+�l��cf�"��u������֨��)�U��߈Ռ���hf����Zf����2��/��<�J��-�e��(�F.�D�O�_�"������S]�@j�L�������wQY���S��Z����pI�WQ�q��}�M�=�ch�zG���%J��2'���x�� U�>0pL�"�#��
��8bο�}v���"R[o\j	[%�9͜O��c|�K�ds}�ٵ'B��7�wA̓�E-�*(���E*\�){�����aŸ�ܳ����H�Fy�׀�!�P.�ȔX�r�%�&�J����Wl'����l�s�Q5�$#i�<�������^�I�}l<�k�@�X2�A:��&�Z� ��e��9��;x��R3�3Oo7����3$�g��@R�<����I~B񗬹Ywu�ׂ���[��JeP�0t
��R ����9Ρ ԃ*��b�gRU����L��L�!l�_�6����T;n!��G
�Gp�{��{�!S��7Y}�~����=���o@��L7�9�]b z1���ևv�`Ȃb ��|�/2kC����/Z#vw��~�U���d3�������}� ��.�W�q����N��1��IS�l�ϟ�9�D��;�EA6]3�g�Ձ�sҋ0=~�<5[����fG97���REL��.zѿt�̣\m�/�\�ē�]o���_�I���hW�
��Jn�S�t=�=Q#�ɔki�dݰ����Wy1��<��۱���|���΂ j�<�7��P	��%W���8�#�o1H������I�e�η���&��
s��o�i����=_�SmL}�������?p�~t���Q�/������kȥɲM���S3�vJ������M�:Y�/��cǫ�=�~f����]|4�V'��(�t��:���{ƹ�@��c�bm�i��<\Wr�9�C�Ч����$M���ń\�+���(�6xA�U�����S��Y/M���P��7 ���b[�	�z����W�5����JN����?
���c/��}zl��	Ϡ�>wZ2⁸��Zb'ȥ �_Y5�ӧB����;�+���_��>�-1�F�5����j�b���F���~���y�d�#����Q���_��an]6���B���Hx�t��B��ㅾ��0�	��1v��d�[����pb�\��J�x�:��{��2[۞`�?M]�.�]����ҙ�&��[g�K�4K�Z��EZ�o�zR��e��9^\�6�MY\�#��o�~Js%�]��ȅe9�3�b�R0��H�_��4T��U?Gv���C��nM�G,���}3h��0��ˮ�t?���`��s96