��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� rā�SZ )����C.��&0C]�-��[�3�-���+��պݣ�k�J�vo`�A�����f����u�X���v�=�а���]Q�Wۿ�߸�=_Q�X����j>��Zw�K��SvX��ƥ.���#�����Z�0���#7{��\S$��@1I�QX~TQ�E��db����۰� ���>0�%�9�j汈��}��1� ��2���h�G��SeY�a���	'<x�p��k�H`�H�j^y�0�s�78+���ֳ�`�R3dW��_��{p[�?$�s0��#�zS�_��bH
�c�p�IL7]� |����Q�� ��Rr���=��E즕2%�����`�^��l�q-�]�p��jf��Ӽ-f%H���ȳ�>��+���M�71��4_�) 3�46h�rb�J�W� k�h~K0�>P$�_n)���5�r�j��W�J&޴o��$>��6��ŀ�;A~<6P��K�~��f��*I
�Z��}`q���ApC��n���g���3��-�іrO�mF���,�$��@�BI�q�}��Ȥ֐����î�䂧��@������U���vU������ �T#K@f�㯁����|95<@���+�-�)�����K���FI�k���*@�m&���
���ma1[�2�u�I�\�U�yu���o�|��2����;�W�W�}P�K>%5�'�8���׫=����k��,�t�M�0�8]q3���N���GvZ�i�+ C�e
��Ќ�S�v<%���q��e_��
�k�夞��>ZO7E~��5k�TW Aod��eE���G���ɑ-'���?�G$����ќ����8ɸ+ 5ʗ���l�d��,�J�
�^�3b,�����J����#n�zK����z�&��;|�\�^���'e�W�����">�w*	FO�Δ��v���I�h���/�*n
�0Zy�����O����z*����2�:�AԶ���U��͆[�Ϣb&�4$56��5Q�=�d�
��
���L��p7�z�Sz�<]�����Q+���%��l;�����pSGީ��}]�u�g:�5ro���+�-䁴��s�9��|�hr�:,��Z�Y��~��oh9�kD�?��I:p� 50��ȞRzѽ�^���	y(qL�z9�y�F�4��d����Y|n�$��[��qC�w�xd�?|�K*3EӇ�}�ή��,��jYʁ��G��(��tE�@a3���MS�(E�?�-fY����^3L�*�A+0�0%l�"����d8��.03�ČE�c>�V�ـí�<�~��L����f*��i<-���ʶ����{��*��A�h'C\����衺��O��zu_W�ޟz�O��� QjyU�� �kqh��O����NM�۴�LZ;H;̾|�p�
� 6��:��ԍpK���n�h��s��2������'�I��sP(v�]�ᮾڀ|�x]�w���%�0'ؤ�d�������xQ��� �p�٨4S<�|�O>�����֚���E�	wa��4��c�x)���Uy�j]k��nFU�ﳋ�-Ѹ��Q�ov��%����駘&�(��K�rן�k��-K�$�9��"�HVb8��=]r�Y)9�.�����J��w�����@��
8��/w���fўX(��"X��"��+�N+���V���>���`��.b��#��! &T$��%D6�C�ؓd	�@������=���<u3&��e6�z�ElT�Ρ��o!Ul?���f<y��3�O����b� ��f`�~�!������g�]|�HiD��8�-��ʁ&�@f5}���,�7�ڔ�V��>{<�v�d:�@O��qKl�.�����7��y<M�������a�+�.F6H�I���S���6Z�vg�	o%��[���%�e���󕎸@��w1��Pn��L�t3غ��'lj�]⪶��BNؽ=��Lt�nU�4�M�C��>�%B�S��\Ku���#l��/'�Y6��V�+�T�f�����B��:=�w�;�:�ǿK����"2˭��G�������pP�y[��Mʱ�q9���zzgd�vPLJn+ ���tK��C����G�<�����=��J��ìBD��ȠjЂ�#��%YW%�>aZ��8���u�mnն�5,����Ke*Ƴ	G���q"X��װ��d���O§[�ɌQfۤ����&�����1@Y�����f����) �*K�C&��cwp�$I��b\��䰸�m<�)�*����l:uE�xu�u;
*�9
ʴ��:��J��K%���?
!N�w�����F�8e���L�G}���ak��7)yܰW�@�������4�B�^��`�;�ʀ��������`�\.UN�D��dCl��H�l��S*[��_oɻ��K�9�YI��(�O�/����cF� ǐ�W`��4��IHWN����pE�E��t�6Y'q/}��9�\�E�vt}'�.�)$H�qb�<l=*0e?����"�\�3+=9���{0/��h���I����
3�0��BW������
Je�1|��Xu�Pu1BB�i���T�=���7��:�����P����6eιH%��s�$$|�:� u�S��߄_�%���M���e�~҈ہ�"0��z�[�8���YP3*�NU8��4����Cj8 �ԗ�?��V�F7�1�}k�4�(a��
G��N�i;Z�Yv��m(���=���/�)���3T�|��j��xOeH�v�Ц�u�����������DB.�޸�g�Drh"�}&�� _�{�=#v9�;i�&
X4u:1g��#0�a��(�\x�>���k�=;�Q%�gg���W'Њz�f ��2��:X�W�����ܽ圩�r��c�Y'w�l�0�E�W'�'aҷ�ɽ�/f��E�;��%�H��j�O��5��X���ٵ`��x�ܦ�M@�w���(���;(��O΢�~l�6f����̲I3��� �{�nf�e7���	k*66�Ng����� ������o��[O_��.u �9��5^�&1㒇�i%t�d2l�=%�2�	p�и|%Ԯ2i�Ļb��@���b�F�q�\��"�Q?�ZK[>��|Zy��ߓ�����<�s�pTP�6�hUZ�����W�(mj���݅�RߠfA��*5	;��oh�^mr%0�4�f��%,�-W�B}:�o(	�uĶP�1��E<n��龛���蟧���܏�u�[a�n2\Ӌ���c�۸t]�����x;��KS��N�j�E�g��R��b�\zE&��j�����ʢ���Z|��Ebr�+yM��=��{�bڊ�R�A4p����Mty�oǩ��Jz<�|��xv�)-������(�'	�Ԉ�u�;�޹�� `Sq%�o]��'+ͥc��]�\jǷ��WX�gP�Z�FSr0��Ƀ�c����(�7U�*�83�j���{�w��܂����L����;\��pFOG'yQ��Q�B�d��#�7`ͤlv1��"d����C=探f�� >Jox؎g^��Gs��	An̰�J�e�PG���z��ޤ/Ap�#:�%^�������8��Gy��7﫤k�����g�,%�m�O��{LJ�^wb8R�R(��$�
�D��(��UM*�s̾��f<�pC҂�+fX6N�
(~�<��G��~X���s�ϴF��G��@(�V� O\�yt'��:����6��#$���S����'
*X���ƽ�.k ����E,�SX�d��`J��?ಷ̉I�_�> ���11�M�%�e�E|WT��9��c�5�G��d:v|e�����0�=~v
	S(�a������H�@�
���$OTS�|$c!����t��v}N|zw'd9��s��F�qc���H�Z�-2��0kab"�oҺ
Z6�?��KYcQ��3\Mk�X�y�_�0Z����~|��K ʎo������@�C���2��w� R��j���}1�s�R�v���i�TV@>�p�������a����Pg"��\�<�s��q�X��D��I�,_�9*���t;Y+�� YB5��1q���4%�!h3�6�b�\4��oY�~���X� b���&7-Z<t��e��=�F�\�2����uZ��<�Q}X�<��0���d`ȮY��0���x�7�/�+�7�(�YJ8�9���n�p����k�Z৅<5a�{�Vx*6�P��L��L���9�ە�F���u�-!D�O�H{�0=J��Ō���X�@񈔑p"�� p��z׋��u��-���j�� ݴ���~��ѱ���#㓬�����9��y�4��vu�Ǎ|��o�8!|kĉ۹X.���nd��B�Zw!%��;ʽཽ���m��E4�� z�x��9�3�b�m�4��opm=+
l�}����&J�T%ѯr��wOˬ�C>
e�SY��~� ���p������6���r�p���DN�R;�)��t'�eJF4W������-��B�t�+&�L��������a�ß?f����A||nW#TDW���8I�x&��{m���5ȹ��\�;��A���&Y�����7ӯ��H�澌��N�z�O\�m�Vpv��ƙ�(��wԜ��+TRC�kk3}��hJ��bB��N1���ӊ��Y�Hqz� Η}p�C+�Ǿ����h.��'ƭs*�D�R���"��>j�{&Y���l��P��s7/�Q����g��N�/\��m`?�ĸj��Ɯ�̯.�f�\����y�z�
����a�0�����F��Y���<�V���_#< �r(���V��lUTV�v�˙Y8����x�o��-#K����u���2���S1�"q&F �M���L�pONL�?�Ȩ~�-���N��-�9Ě�w�C�P�,Y��`�T��vtĢ���N�P!ʭ������p�nv��M�M��i$:?��\T���²�F�j�;G�g�&��v�y#�F�?�ǔ��cjoc���C�h%!�<)�l�e��4����f-�U�v�m׳�Y=]I� �) �p=.΄V�n�o�U��o됰:u.���V�D��號0�<8��R�����H�_�����lm��~<���]H�c5�
��Z�����t�8^���6��jL��:V�v��3O���d����#�\.�vEq%@AfiW
^���Г�Hz	���Ǎg��x/5+��6i5$x�e�})�����>��~rQ��=����5[֤&<a ��\� $���//�#�.��y�(�1��q����m=\?�ȭ�� ����E%����4�H���a��T�J����k�[.M26�`�IE(������I���[c�b��BpR��p�Z�-����I�i��%:��&��ъ�s��EY�r��@3	�o��pv8ؓ����	;�O2�
c;'�1�����6��^2?��lQC)eH�G|ى]o�J��5-Zmy���s^ߠ�'��Ĕ-�y�B�*h^n�������X]��}>�5<�_����w������jX>d;>�E�A~Zhs:I�Q��Af$<��	;ѵ"�������VV��F��D���6$�3�E+��E���3��ϋ�'�e�OCt��[䲒e�B��ȸ����|7���sߠe�Lh�<������+KeCQK�ƩH�U��� s��!�X]�N\E��)��r�^x'm�Z5�b*�O�>�via�C�\Re�ʖ���2��xa,4�"��v��^��e�_l�s91�T��AW��K@�¼h�>��`��P��ƶ�6âu����?3�!�_H ��������ag��]y�Z�}��
��Ҝ�l5x�8�q�	4#9��Y&Pqy�s�0��Z��7�@�f£/Η�%�5����II`�,�b���n�}���$Il���+���I�&��8�`<'������%�{3x��lHk�6��[�Tc�[j xd����^�_���c� �FY����kL��ϱ�/��BƑ��~>�s0d�j��x;jh����K^T��g*a��6��]���ߵ "t�h-3
��]�/>W?:����z'J��ZQc,}ժ���c��R,����~���i�{뎳�q+�57�����<C�I�3"xG��Z��<C,3(�S�Dn�eY��ܻ�-��/o{eд�-��w��t+?�k$�(>:�fy�|��N��4(Zv��|�W�����.Iw��-�-A����j�XK��._D�Ly+��f �	��/���`j�4�Yj�s2�p����̯�Z�@�jA���\F=?�og1� ��ے_��3���+�迾��N+���I[W�F��k�g����@�U��۬5:��j��S6&?�u�)}��ɽK��'ˢ=�	`(%��u��L������h��6L�2�"4���<��>n�y8�"H��	
�	]�L�A|Ҋӆ	��!� A���Gďch�h�b�Ue��u�T{D^��H�TM��� 
����6�3�g�P��A�)"MA��:�v�Ĝ~)�8җyyԱV�����4[�s�XY��:��R~#W���DT;p��1�-���X���n� �cն>0�_x�;��7������E��#��`���>�˩Ji�4S��r�ca�t���R�o�ހ�=���܂�Ò:��3�����	9�wA�%�bX���N%!l!Fx9&�aQ���[���na�΂��'���'Dt*�e�������B9Q~\�OT�3A�%oi��F�q~�qN�bm��(��N�bp��Bಐ�"J�[��k��H2�.^���9���y�ϳ�o��\aD6F$��!LZ��4y�^j�.�ճ�eʸ�ҿ�lQs?'���ɟ5��{GS\ �%�h}��g{�&�.��J>�ӕ8������,��r����8$	t�X�1İ�V*l���$��������Tz�>fzR(G`��.H(��' �X�J�䅖��G4��
4��nc�x
�����B�D9�M����WH��<q�;L�Mz``�s�h�a��C����?4����jȐn��Qn��l>�O�YH���z<Jo.�s�^�O͟�E��@EqX�!'��J��V5k�<���uŇ"%i�쬷�4��YHѸ��
M�W���jH�� @�ӸfΓS�����̆��o��W�����1y��\�Vx=䕯�[��<��j�	��~��S60���q�Q=3G�$�xyRS��������޶��`ɗͯ��UN�.�"�,��Æh�Ylc�����>��>�I��R��R�_Ks�E��`��Q���.�]̪��S�C~�����
�8��F�(p�)�Q7�z��UT�ѐS�.z�������t=,����J�$���ả����7K��t��2�cm��s�΋��2���d�f<�_C�`]o����;�
}wv����l�=t/�t������X�52]��.Cܩ'F����I�EWH��g�]Z4jX��Ebc�E	bڴ�^{j����{��>S:��=c>k�+&������Jznج��!���܄?�$�WP���B_�k�0xT�P{l?b���醜�H��ظ⦎a��+�/�cu��H�����Љמ�5��n"v�^q��L�Nޑ���,�����!.�naU���-�WR�cu�-�U��fJ��En�����'5؋31B2�Ģ�d �� ��݂�;z�������������]�$"���M����=��C�#Q�I�'�M��ɧ�Vm{�o�a/�@�(;+�~�%���Zr	��P&��>��p>~D��?��+�+B0�p����'G�i� �t����Z�� ���<��������Q?z�����ݑ��ZB�1ƿ�͖ք��Q߻�R�����V�R������X����_�d�8���OxH�>�5ig��VJK�S�@(y"K����[����V�q����W����Q|���;8�/K�<�"������z�ɕ�v�>Zle���8�H3d��O���A��T�QȊ���҅<	��P�p���Ӿ0�׆���g�
�Yw��� ���⁆��o�)��R�/���)�F7�	Rŗ�〲<�ܰ5���{���m`rp�͖�����Sc@7aj;ٰy����<.Y��͵��-.�cX��c��Ù�]���'Se�xX�R凴r[���p�@�����a"��O}l�k�^�������l/0���4^<��Ǝ������f��ٛ{o\��_���(�0T�qAOM��X <���B2�ѕ����Ӎ�T� 
%�9��l1P�x�9��L�@NcR];����
������+�%�3��j��+ڠ��iۡt�5��F)���꥜�Բ���\���I��Zli,��qy+Oܸ��@�z���k����Q4:�?h�?J�n�&�v�v˄�S����e���`nA�|O4n?�݉+�ϭ�IqǓ���{���zQ�;K�X����7Q@_Ghh�R�3cj5�ks��3$��-�-�d�����?>�SWH��D��/%Q��Q�YfJ�L�Q7��6}`�m����B��*�`g ʅ�y(�0k���;�-���5��r�\-�Kv � نӴj���Y�3_��?ЯC~�%[2����	���Ȫ���@"&�Z�QV)/�p����'Gl\��f(r����4�ާwk�-Q�҄�p#dK�9Ȟ�Rjh�l7���`�K����i�y��/P��Lh߂��8����{nh�nO��,���D�u�E.�͊�o�3�4�����8���j��lYS�]l�4��.��A�KE�$In<��=߶�a��6f�;���lq��QDx�\)OOm���@8§������&!.SbB��������(�tf-�p� ��^v���:S��yt8�%Tc���z��Ϩ�f̨HW�~�;���y��E�J��*�_ƃ�5�'r�
�����h�$p�d��_��@@�cሇP�CS�ӆ��PA���q8`�Cj�yD���^f .	X.����n���yݗ���̵!��L��ǎ�_�|����m:!�C1g^��������NY�Kn�h����*�/�ۧ����w��of���P�x�J7l����9���o-u���|m��f,��L�4���0�t{oٻ�4T�Q_�~�G)��8��ȷ�;��iD��û���S�p�T��1�٫y�3���M��w���oa��
܇Qg���-���h�)]��u�ǒOt������ῶ�Db��y�]^��7T�������:GЃi�	c�����F"��m����ծ�4?*�F��a�nb��B���$��i9^��r�O�L(�{���g�)��K�"��\��ZgVv9�O1W�edL�0���>m�kXc�7�C�wa�s�3P�=P�Xe��Q�����+��Z�ͥbS{:����~%����zOT��z� mFI �j��Ԙ�E��2����ٜh�����XFt���h+��}Q��0��,��Eڈsn'����致���y�ם!�b���D��z��]MT��0	>����ν��e�'����R)�
\�0/՚�����B�u�}���~���e�	����7Ms���G4�X��kQ�G2�iwfm6C`�5��
1�<�P�$��i�/�+N %e.܊QP�#'��b2��e�%����D�9cYrW�1Y�`��JXȫ���d�Q�+o���y�H�C�M�֌Dq��})�N{�"��8�F���r+�P����?�4(LC۞i��̓�`x�?�������Z�k\9�:��NO���{�6k2c��h�X(�;H`F1C?+Z^��<�,*�{T6J��E��f��g#!L�83�F_&��	^�;�H
��+�@\���?����3V�n�X@�d�)BZ�F�W�f��0�'�B:����:3��N쪄N}0#&+�&AE���k38`S��҃Ëe�c�q-�$�}����>4`lx����?&
���`����R~}���C�>����e����:��{̥^�:�IK�l��u�?�!�&;,X�Wc�M��
������{|,�M<2�N�zP�H�s�u����3�.��`e��(]���n��J����8�3��R�tn�-m�y=����b��a��L?��*e-���Ť��N��:4p�̫|��sG��,���Bg�e����*L���,@���-�?������Qqk8��]{��p��[��GݛH�<<��@Xd��,gt�e�'�'͋�Sa���ᒜ��*d��E`s}����a�$W�Jx&��~�����H��t��$��$���
E��I�̈́�`�n�>
~ c�N�'�p<��[�6���wM58
X��cr�
2�\F�3Z�-�7�i^:{%VG:��aĊ�_��[G���w�������G�?3�[�1�U�cԨ�<��%�Gp��q��g���(�d��O����/DgRt?]8��A��#��(ΰ/��Y%�~"<P{�.)�'(�U_P�%i�^f����x�mKT���bdn��~���7an�H�+ӕ2|f�-�QLܙ��^�w�ҨB��w�Z�h�di3q)*=	�b���F� �#]�쎢Y�"jWx�.Dl�;n���٠�Җ�74�fμG�*�uo}@(�l�$��)����r�2ߤF<[FsS$sf>��9�+ɮ�E�%]�oS�Pg#��פ__bh�Ͻ �ߓ:}P�R��@�T�M�s	s��٣h��n�m�3�BkZE��
�x��j�
���s��V9��'"84��uD ���o�nS(���_����)g��S�  ��wS1��~$׻�C��G��jKٿ����tp$��Ɂ���؛7c�(N�#��Q;qD�~�F�� I���K�B�7;��()�]}�E�z}�c����|u����/5��a�n�'0��֝v�[*e ����jS�3JZ�գ,G�yAB5!Z�D�>��s���π>"m��0rY�Y��UՑ;r	�ƀF�ҥ� �����?߉�)�M��W�mY�H�F�X��_��<r=��/�ڈ��~*��Zw�j%�j먰MQ% C��'�Y3Y�@��~�L\��f\��6�t�g��"Cr��\��~mk������V�#͹�Չ�)h�b�'-���/&��'��K�3��(n�N�Á��(
E�b�x�kD��ŕ}�ܺ�a�y,eM^�2ك�G1�:J_Pk���W�WV����M�r���*8�8*g�ǿ�X�h
|�݉E�
��V_mN*�aGOkO;����S��?7� mj}��*����t��o�v�b�A�7��F������jKN���@Vq�.��B$��̳��S��G�
U������]��a=�Y�7	�Ԉ�k������Y`j;傞:�G�N`xH��/�d@��HR���%�w�wt�(ki�96i���� �X!��+�I�J�GS�Z��j�P���,�Z��zaK���<��9\/�Y&��ɚIn�hT�&į���s��t��C� U���yG��L�t4�̸��s%;�H���a��]9��
�2�M��<l�	���_�U�;�Osx!�Ru��s���Y��e��O�}��x�Z����KX\dP�ѽ\2☟� ��hYX:���m��vD�i�DZLI��v(pp)j���v^IU��򓺲�qݗ��^���/�`��g'X�2d�ʷo�vG�`��id6Y1�%�ƍ:�d��蒵`:�7�G�S��'M���ĩ���os�ܐl���		���x��`��*R��#��F�0&�}DǴ^y<,4H�a�w� �Kzkn���ZZ�r��/7�����C�z|��'`�;;�}�f(����?Bǰ�_~Y�����e���\~ :���s� ڤl�>qE�B��csX0$�P o�[Ǻ�=��pه����֌�@}��E�Ī/���i�ޠ��}�p�x�e�ޜ}l�_*�V���.�ݔ��z�~� P�K�\��?&�F��4 n���(�"��?&1��۲����5�_dv�e8����*_���<T��v�&!0ǃ�O��1g��A���닺��W�bEs�O���dA�|[TL�xQ$҂hįY� �,=�Yl*~V-m��Rh�g�V�J��RLȼ,g��0����ӵ�rV��Ŝ�1��q*	��U��#���Wቴa��<���w0H,�~�R<JC>�z���S�'��9)>�c�6��EHmm�ֲb��;�����{���v�����"ٖ)�@�(�"���y�<��۳��v�t�Q��#im,,�Y��-?�V�w������<��d�|���9�6pk1=�p�酓�j��f��x,Đ�0p��%��`R/�#{��y��?���*fG��!��o���z
]����_}���f7_�B�nG�*�S�2 e�<)t�]��3�������h{*D��\���7N�Tʤc(���xЕwB'd�%n��ȃ���=���y�Z7�(�k��Nt���S/��L��7j@�D:1�*ɀhUt?QU��g5M���gs�R�T�j_�Y����s��/5����9�^>i�_�,�3��u�����S\�e�O�|n��4V���:�A컪�Rq���s�,'˳z�QN'W��j�HO~�7�b<��]$4Y�4i��bg������ꘀ3[Yη�
����E�X!��W��#�M�(e����	�����v��p�7~�	�d�6�����c=�ɸzB�bz�l�¨G���dV�Ӝ;��c4��_3L�c��?т+�q�Q���z~�_��	܍����r�M��k�s��S�#�=���Op�>:���
rc�AZ;r3��5�h�����[��(��]$M�Mpj[guSC&)�8�/�Կ u�m�y٭�[1T�1�J��W�����4|��_��-�M����ʯBr�r�6^
h���qW����jZ��7}q�������i��v��������~�'{���p?�,�9��"N5Y8�n*��� Zm"Pa���T*�\��D�䶶���d*�}��� ��wnp��s�JW��[bv�.RKWњyױ�0eh��(P��vw6����oy&�2���A+@A������;��h?P�)�ہ���t����5�]��Y�{�����Sk���Lg�V��1�����W��U`���z���9�S	�$���|Q=\5i�iiWh��hS?X��Z��`Мy���&Gp-����!��[�"�"�rK�Ĝ�ۚ�'���&�1!����`Y��D%D�ԃ?��� 8X.b��yK��`��+NqE�[�*��y9��YW�r	�	?�+/)E>���Ԯc�%����h��������X6��+�AH�ˤ;'�4��1ST���Z*.������4D5��(����h��,zF�S��z��-��>Y��}(?����]�O ����r�@�Z5�dݘSA���[��>3���)��p�Q:!g3�+�ߛt�np5:����v gC�����*5wDҾ��)�=0CV�U�LMvs��M�k
�.���姇��._�c���)���
NX�Y�<� b�r�5���u���-'���W�W�Њ����u�a"��r�g$ucI�k5����!֟�[\�:�0��04R��[A��@u��(YR����0�姅��'�u��4B�Ͻ�ո�T
6��#�!�u���t� �?����N�N=A܆v��;��AC�u��2��4hڑ��� ��w�~����f6��d��3��')BLb��aw8%yЅ�HA�����ۋӈ�^�	|0תϚXb���E���ǹ�Ŋ�£��GE)p���*~,�sV���N�54�=|~��a%�@D?���AN&�������eʁ	=�34�y'��
p�7C�2�͡��9Ȧ�ݾFfiO�����%`pArrj����{�(���6��-&T_�Vn�x��S��m1�$��0��&D=i7vo�+��$Hs����2]X�!��#�vs<5��U�)��'7���phQ��fqY�7/�*���Rj�h��?��~Eu����Yb>ס4*��OR��􆢃){ ���ar�ܛ�J���L��L�B��!0�Z^g�1j��TqO���q&�K���R50��܈��r���B��;��^º�V�`��q�"��0�����S�Me���J �Ty�"���+�S�K�����M���~�28�G����AR�1z�)��+gP�������^��L��2�f�Q���aS����v�4n�z)����"9��y�0`��W��\����)Z!�n�w��ߢ���[�ң�-{h��S�j.���(��
�h�Git����Z�r�'��#ϔ>���>��ǉ ��J��cl�~�1��G���l^6N�`�քYχ�DM֛��r��Sp��?SQ������� �-�I/�d�U���u�DM�������~Gp7��!�/�T ��2��=[>$�$���a:};�<7߈z��@�C�J�����M����3Q��l
��`�3Qc��cJ ʞZ��Ğ^�(G:؇P���{5}i��.�DA�qt����7��-Sd����f�,�_�f���B���p���sL^�S-�xF�`ʲ)�{���4��� b����.ȱ��Q��28ϻ�������Jޥ��� ������si�/�2����_ L�<=��^#0�j� �8���ĒY����� e�m��\�=��9Aڔ�O
�q+O�0��>q�ߣ=}���.-�Qs������MKɍ��H'�2:������i�׽�a��V�g�?����#�9L���K�`l�a�rR� 4�O����x.2�T�����N�e��J&3/���2�����۰��� >��dIʼĪ�2��R?�^7G�N�gs{oY}�;�/$����x����s�`���U�r�_�i=�"�����X�����b�S�K^�=���A$� &���'� 4���t��h[�3�r���=��7;;vg�����.7����p�|!���)S�7��4��д�]���Ǐ��P�6�Ē�p�{# ���ۤف���v;����{{ܼ��cu�[5�H� A�T�~X�C�T&ߴb\9�>������A5)=L>���s��-~i���t�73��<���U���Hϐ��Wc��ze
��������)��V|�C^gq>
>R�&��!s`�_�����G��EI>'y���:?�� �&�*t%���f�ߒ�����6A��A/
�|�)E�[<bEp��G�gy�rY��N��H��x6�o/\��'J���6;�P�v�bH���lvq0�U
���9�4�כe�l	[�Oƃ9O�&�ݯu>�#������$�`gyn���r.��	}�/�qL�W$�j��`2MK�BZP��[[��XJ�q�Ӱ����(�hȥpbG��� ��%�'��OK���o����q�>''���Cz�@��,��S�0����)��\1�����Mm��}�"4?��K:�Q&%�����(e��EI6���Ui
�rJ\�l���?Ѓ�R��D�Vc�� @E��4p5���w�%�U0�����n�lLK[=�Q#��u3�(��MM+`�����r S$6������c����3�1�^�G�_��07��W(yn-iqF�ϙ��<k����n�U2O`�-���D���%_8fYA�؂�����C������.<Bu�N��U8���,�c���w��P��L��fd�D$��U����c��^�����c�IT�f�����*d���b���;�N��h��уYxW�.g�#^R�E����S�"�X�<%Z�)��V�}L �:d��{�pγ��"�;(,�����3����{-�J�_)��Mm���ֳ̜�mLP�l����	ubD�;��02]�B?�d��yx�D�0����(�Ϋ�Ei��y�e��u�({���V4�*��
�2�P�_��` 7ܤɶ<`'�B"}�TFi�z���G� i� �LOAi�B ��
Q�)����|�HZ�!9b"����,������,�*�<*�p���?�<ǒz�O�C���r/������*��}MIw�	Mk�L�웉��i��]�ǽ�L.R��q���ۼ5�P��	*�b�PT����ޣ?�!tS��齃 �&@b��PT�1��i�iƴ�	�<0��8��2�xYm�ruU�9����?*�u���e��C��[�wBɘ�nuG�F�Ǩ�<��N��E}.�7�����A��(����j�"+��۝�G���<3��ʞ��2�= �:4�]gW]ޢr	�3�n6��ۑj;�sU���
�8�m�����	+�f;#I[!���5�ר�����6p����$7���b��>�L^C�]��Kr�>F��7��C��vN�*#A~��6���3
|�m��P�<wz������`7\�s��~�3�Ꮥ�5���s���B�S�e��F���[���@�)�%co���ؿ>&��d�s��f�ą�j�%v ���'H��y�]�G�"�صKb}')����ez��@�r������s���=�w��fu�p'eJ��F��i��U]v�a�!�m���pZ��x�Iʜ�����y�.S\����h��ߖ��� %�P�f[0YO]�Q?��r��r(�L랲H赬���9˛�w�wK����	>�>��S�����&�w�Y��#��ԱP�w�ÀB�U:-~bh��~kIY����}�,h�����9�X��M-m���"�W�������KK�d3wg�8FYh\k�Fo�u�O���� ����$
����u��؇<)!t�A��t45E:'�R���b�N��6�N�ɔ�|��E��w=���$x̍�d���7 ҩ���?�s�ZA`���ʳn�m� �bJ���|�6^8O��Y�s��Q(n��qHd[�p���?ݔ�"P�iժ"��j�L)n����2-�	�@��t�	�����Z����f�%��2���4=tK-8�r��d�Yv�X]?��(�(,��u)�-|���E�u����l�g�I�
r�e:h����c�dCwt�xe�{b.�_A\t��d�A3��G�����g�����gǘv^p��g�.�W��������Z1�a�|)w_e�s��|��A���s���X��eCb�60<��i�嘥7rt���������",'�\��#(M�� cuJ���h���,�;Wh�y~�=�!x�YQ2����Olf	�s��/��YD^���i9��4f�WR��*� ��}*���dy���wXҚ�L*Ϥ]�V�'AO�v��T�+�G�+�ˮ�M�\-����!㑽{n��K+��X�4C��%��1	�9�~$�=�ZO.���B����/��,!qC���K�$j%�UQK�CΒ�*�ǩ�5e
��q�jxu���ѽe\V��4�j����Y���u4��}�ax��v��>�ֽ��Z+h�r$��-�*9�VP�7�����(������}4��p�?�#��s��L����D�	o�? �n1m��t�L ��������(P�S�d��9Ro$�A?�<cM}�(/���a��� ��{m܅����� �1�F-v3���(p
`�s���|�1b���n��Пդ�;� �V�kͧ����h<���ù��a|��]��p��}���e%ݨ^L�h����q.YDB���)��V0:�D�X����f���U���[���lV�L��%��������x�R��?�g3�P�n�"ar[�L�u�B*�������Io����^�p��Y�#b�U�'{��H�G�
V^y�����$�%�f�u���O?;J�Uj��&�sT���o|g��c��gl.B�y=����-v/k˫���T,z�%���j� ��0:��]w�&(�����z�\�f�L��C��N$��$j�ʐe�b|���T�E%|�A29��U���ٙ���8 ���?hk���j�/(%u95���jF��Q)��@׹]�ֽ����q��ϲ�|�_)��ޚ�5	�� ���l�\��5�x�nb�dz�s�)`DG��t"蟩)3 ��w����x��E��sc�ZY���2�|] {�u�`�A�h�r*�ؔ�+{��E(��n� ��
���R}�MW_����"�{�3���u7w�m�~�vgN(a��� �2����S#bO&���j@��]`���
�R3�__��Һ4�4��`�������ߝ*�
��������<&��\]�[3'7��Fy��y�l
��K1C�L��%@}���������ȄGv	�h��������i3|�mȂ� ��/��,9�L8��
T�ok)�~��2"Y�,
�H
����8ҖZ��SX�v�)��t��
Pa8[@��`*�)ɀlI;;��Ǘ'TZ
K`����\�k_��F3�bc�/�"%"&�<<�x�f�w���a�n�v�k��s9OAKi�i%�x)C�0l5>��s0�u�03.V,�~��\�nQ���"5:�γ�m�_K�y��<=��F�'gH��*�\���T.9��"�e����x�XA-Q�Jʕ���D�Q��XАm<��Jy3
������MP�ɘb2���M�]�l "f�U���eW�ul�j�q�v
�>h��$��aƸfK3�T�<`U���㝊��]�_�42�?�1�,� 틪�S�����҅x�vc,��xstdNm�*�i�:/��Q�{���|B�؊�����_�@˴��0��!��c�BP^�m�2�;>��{m�2^��"k����3�t-S��_��Ȅ�:�o�B%�ag�	��ǆ�TaR^�>�qf�K$����L,L����y���WŇ,2;�r�i��ԠV�J��/p�^2�_��W�8��=;S�PY�Yg��c#-o)��+���� NM��/y a�4`]�'�
�~_�|�M�8)��cm�RE�da�t�eW��tʩ�1WS���~��k�P	-i!����;�g�!E����Ƞ��Yg��X.���X�\�b����CMy���C@�R�#��F@*݅��O���K'6�9I����MA2t���Eۓ|�x�O��1:	�O��B��|��]X&7cO�Q�҇����Fz�������jT)B������S��\Y���
2�5��"w�Q���U�	Ҽ=H;�R�Q8�i���Xy������s`��u�LY�GdjJ@�X���~�.W}\B����{��Ϡ�)��;���WÔ\�A�@	��/<��G���Z��0Y�#)�j�����5�/��g}��$8�܌U!q���R� ��(�';F�:=ӗ�d[���&�@���]��HG�V�a���Ǟ�=�a}a�����I���M
5N��j2��A��C�X|�U-��Di:`.�m��W�Q-�R��wܙbI"'?��O��Ĭ��D]�"���N���AP�IP村m����utkK�u��;6��K?�=��WL ���v�PT|�'Y#�g�nbI����мz\�I9]e����P�L���<���~'���4Mw}Wٴ��ׁ��r��|�!�Oc����,e(v­�o.5����:�Qs�T�Kk��b��Q�s��j��O�Z�HXy]q���sű��2�g��[�Գ�_T��`[[(�Lq	tIGK���t��U���֍����?s���b��5���s7�����ܸ���큶���L��pU&�&):^TO	"�E@����#�O����!�����%��)�U���+�#�6Tu0J�d��`��J��#��>���Ƙ�&�d�O%1L��t+m��?���ؖf�Ϡ��o�u�/9}Ik
��dbR(�1q��V~�u`{T��*��c����)�\�(w�~fm�3D�b�1��!��ߍ^���e�<�H\��q@�]����4�a��m�Z����D�f�K�F�>b}&�-[���#P��熧�U1E��)������!�]�|e��&� �!���T[���@�b�=�B��H��b��Ԣ��P>M�p�|�;&a�N˟Ln�k�K}�*0_;�Mϊi1�!;�F����a���3�B@6�F]�w��M���\���n���GuǷ�}�1��3]RsN���d4�lTc��㤋XK<k��
��!J�{0��
 �jH{'̔��p��ٮO���hӑtfҳ�ċ!���
"km�94:���ʪ��	P��JNq�������~�(�~�q��V���*\�G��aS'�Bؿ�c�GZ�����A� Ja:{��WP�e��k�����c��c2�&�� V9�;�E���۟����d�q�6�p�Tv�Tz������O�Z`��l}_i0Ǖ%?����dT9��[�M�oZv!g��*��k��|�*rL�=g2�n�� ���V@y��Zl.+���O�\1˂Q-�ڡ}
���ͪ�`jʖ�3F��s�~Ѧ�"g��H|�l�.�Xx�FWP�	�(�[k2,K��Zx ׌��H�]�|�d�ho`ǓI �p��e�-�į"f�\���l�a����,%Ca����,dZ��1C6�˼-�6�Vf9�;����{�/�����i�0�dMIr�}�=E����#OnFm�!��J]K+C�hN�=�nB�S(/��!��D����9��ZTq$�o#�㽐�
wXNpPh��sJ�x粹*�Ht���T:�W���jQ�q���9g���EH ��o��,l��n#5�_竟D�0�5�Z|���EV�ב�UE�}V3��Dٷ�޿������ۘ]8_��'B	��I���m��Tw��9��h4TkRA���j����ff/G�b<�At��ʂ�7Ϣ	]���O8T�y���rf,��vbL�d��a�zGT�*���H��!`���)+����>,�ƅ�)��v6�MЌ-L��i�#}ۼ�a�)���<E�6u
F6߆e��LD�hh��P�۶�)�t�2��ͩ�(7��}�-��$ �4V��	���Z�%��G��,44�HN�F�����*���0ǚ5'N��!�rf�\��s�� ԺQ��.��(�X��Ř�aU�gqH���2�8��@1��oi���_g��l)���:��N���F��:�2��������)r��}uŉ)�Ε1�>54B�~�5N=�H��\�.�fM��f��eqȮO-��	�s�8�*m��˻�)�I��WA��f�],���!W��E-b>})����:���v~v��ɯ��[rA��`�^�z)��W-�Kv�@�V�$��i'(@2��\'�B�U��;j����+Li�:W�{�;5hY��W_��T�zw	~ .C��,�0���0��^���#�0z[��s�a�IEd��`	�ڼH��SJx�JL׮pW����Qu��^��&d �C�����K�F���_�sG�� foKp0W��v9(�@Cn�������c"뒔���ITv�f��v�a�'�A��}$)�N��,�ԞeS�_�yc��(P�Xxs����07��]We�J!F�ώ��x8L���y^h\�=T1ź�u8�g��4�>!T2�'�-�N`�B���)a!諅��ـN�7�����~���LM���J��A��l�$M]&bs&Ih�����&�9*HC4������2��.r��"BE���'��x��o�,ɉ.ks5Ԙ$9E���(��`�$E���m&�� �4�"�"j�C�?�)�0|���l���ۭ��$K�,B��`��M����Hiϻ�����C�����Ty���5BӐ�LK�t�%�jm�%�c��@��<!�˩�!B�0��4׻����G�+�rb�w1Z�0�.�9,��}�MX�fΘ@�O�|�RE6�P	�?��9�s��������z^M�ӵ\F"L�
���+��^̫|
�	-*�$��>c`[+pBNٳ����mj�p�A/�/č&.䘍oHͶ��`MZa�P��?���q��j,�>.��m����K�S6t�`i��P�Z���i�7�v�o�m8�\���sè*D���'"��Է;���)5g��nڑʙ�0EV'�~���a3��"���(���9(a����.�?����
{��sĢ ���=�;����vm���Q�X�5Nnx"�����,L����d0w�'�) WHEE
��%H��:Yy�b�*\�.�]ir@����U�	��<�c x�߫�\���=V1u>[� ��r���*3q�ܦt1r�nM�Z�p�u�]�q��}J<�u�:ے��Hŷ�f'�b��t5�*�*�p4�$�e�*Z�G�����#'���A&훲1�{�XY��9T���.X�#��J��2卟���[<��p�i�1޺��%�-ma�dޮ\[�ٳ�F{�1v���iQ�)��	k�\��̈ɴ�!�ݏ�W�=��u	���J�2S��lctBn~�|�UcX�jh�[@Q�<'=�����)>�?9�8ӹ���Uz�PV%���\��oɏ��4�13h�*��ʚ�<�c��f�l0��b��N��n�AR�oF� �0�֧���a��M��3 �`$;a�i!��;8�=�D��4�O����c��;o�����||�w�0�+���/TŒώ�%�K�M;�m�*&��G
�l?�݀�l��F��J�""�E���i���a��!�@0�g:x�Z����ee��H%�hd���=�V�^�2dc�ޠ�B��r~�^bY����
����g���1Mu�V|�G�&t��g�eߌ��a�mؘx�Q����5������#���/S޵�Vַ�;��|��X?�i�1|-���|�K�7�ĥ�p���P�k��sz���Bt+)�u�w��*�wύ> s��f�>-�~Ѡ����@�?S�п�K>@��H=cpEK��5���]1 �sCJ[�K�ԟ��~�Ϗ�@��ٲN
*����O�Წ	�	�HrP[9���v�~�7��(D`k)��f���"�َ�WX�I���1���j"����}"v|@�S�>�0es�)��"Ԗ�C�
P��eY�|Je(�N��1��:���>��c2�*�I���3�uG�@��"��!1��b�Bm�f��}w�c��O܊F<B�f��J����3LF�`Yg\�o���G��12C���>�+�%���9=ף�\�k�[Ex�P�:*6q���-*���8��fY�(�*�F��Z$��8���URt�����ÒV�;e81�#���#�V��J|��d�����U?����ؙ7涏�����1>݈(f�m\��x\�w��)_7���#jq]�ȍ��bu��)M{%���
§�u��b<��i�P�3.�Z�1{��[6G�ug�q(`��KE�7�gh�g�˵噷`
���B�����	F^�oM������1�E.�T��	]y#@L*��>\�ǜ��O�i&�t(����ۢ5�FK�9Q}�M�@�����9,	F��Mz��ha�[2"M���,!>������P@�N����o�.V�ҫO�&������N��c�WpNL���#�]ΒW[�������zY���ygG�.���;M�m�1�H�n?c���rc�L~�K�N2��^�Ū ���s�}�V��ʀ4�^u4�k����׌�&ghF佣O,�V8@�zfK���3��^�������DV��Q��XR_@�ٮz>�(28>��|�3���%%���?~�QPA���]�Tˎ�8I]g4��0�Ɩk^�8,���[���	��MqLJ�-(�=K���8T�*_�?�x�H��l��\���Ba��0�mS�sI�?�zo1�h��@��i2`1������N�@j->qv��s����&�
ܰl~��#�n�c�-���g��rְ����+X+b�>,���Z|�A@;��b�;b�9��c��^wX����ƀ$ �YƩ����Kb_e�PP(�Gj�%��s{;>J�!�%C�*�~j^�%I������}����x�.�b�$\ ȑ��e��P�Gݼ�3��l��J�͟Hi	�@��� �p�ͷ�--R��F�������ٴ	�ʹ*FˈI��?�20�NTzx<t���� �J��;l�7���Wb��C���7/���?�4���u�W��d��;x�\?�y���z	$�