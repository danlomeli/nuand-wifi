��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� rā�SZ )����C.��&0C]�-��[�3�-���+��պݣ�k�J�vo`�A�����f����u�X���v�=�а���]Q�Wۿ�߸�=_Q�X����j>��Zw�K��SvX��ƥ.���#�����Z�0���#7{��\S$��@1I�QX~TQ�E��db����۰� ���>0�%�9�j汈��}��1� ��2���h�G��SeY�a���	'<x�p��k�H`�H�j^y�0�s�78+���ֳ�`�R3dW��_��{p[�?$�s0��#�zS�_��bH
�c�p�IL7]� |����Q�� ��Rr���=��E즕2%�����`�^��l�q-�]�p��jf��Ӽ-f%H���ȳ�>��+���M�71��4_�) 3�46h�rb�J�W� k�h~K0�>P$�_n)���5�r�j��W�J&޴o��$>��6��ŀ�;A~<6P��K�~��f��*I
�Z��}`q���ApC��n���g���3��-�іrO�mF���,�$��@�BI�q�}��Ȥ֐����î�䂧��@������U���vU������ �T#K@f�㯁����|95<@���+�-�)�����K���FI�k���*@�m&���
���ma1[�2�u�I�\�U�yu���o�|��2����;�W�W�}P�K>%5�'�8���׫=����k��,�t�M�0�8]q3���N���GvZ�#z�HM���5[mWJ�S��1	����,8�5 -�3b+�ꎖ�jiy���(��[�8��a��:��c�j␐|���$��O��5�k=�-|��GG妄6��TzO.�4�,��OJn�9��߶�p�+��0���o���&�(j$�����x�f��o	S�n��/���+~&(~b<"bW7��^a�t�7J�;����=����o>k�UnO�NU�j4� .����wK� �G�딋d��Y2O50����U�^7���X�`�]�'�v�f�a�:�&y`��uFft�B�����ٕ�gR�� ��M��?��T�s�N�ۗ����=���R�(�����9��gLk2H'b��L�Z:��JG�2�1���Ak�V�B��6o�p�8�࢒�F�3��	�����}��F=�h��M��5�VO�7j��9 ��QR�0�ᦸ�\���L�n���;�����4���߇�̛��Y�X<���R8#PD���������}��$�F����AH��Z�/���"D��~c��gc�"��H}��/G�]m��v���kƖ�$��2+>��Nf�P��$Kgum'wJy��G��lhK��� f<�:�&��	G��mp�ͫ�^����i�B�EA"�����`�xL�� "���+�7�$��-�HÁ�b��3h�����V��2n���qFN0��� }�̄����}��INL}[�#㽋С���W�@�=����2��8�ޜ %�{��V=uQU���R��g'�q k3���,���O�ԕb��/���mL�iʅ#���G\�?-�W%M�-!�{�~~k�*�.`��Q6%�06Z�5��t�֓�A�T�ɋ����`0�P���i%u�M{�V״����2ceZM�0{�L*"W���Oe2-���Rh1�p[�`C2�MS�-ڛO&�,%�i�^����7A�Hn�̡�(�gP��c������ۂ`���4v0�T�on���i_8�3�ǂ�	Cư�g}�4��ph^F�M�{�( #�TK4v8"��z8���77�^6����2�ܧaE��
�n�C}۫x�p��;L�V
�h��c!Ozh�R����T��+l\#Tg�	�0E啚n+�B'��3�A�a�F�X#a��-T�i�H5Ǆݰ⻟�|6[L�wD{W�V$�k܌��:��@���ΰcS2j�,hL�C�ɝU�3L`�치�ӌ3Ʋ�e�G�	�^��??ԭ���Y�`Q���2(v�L�J {)��%�w6��D'�Y#���-�2&m�'1@�q� �Tz���ӡ,hM��y��wv{�U�e��� ����d���2��!,�ӑ Z&��K�%�;�W����ZdQ�����#:mG~Wr��8q�]�h�wf"���38�{�I4:�'5����,��\|��E�4V��&�
LtA/4��r������O�IG����6�D�.�����=�1��sU� �Ȱ;V��P�J��y�Hæ=�Y��Tb �b.���`�w��r/G/�l1�!��r/g���ڽ���y�J �.��:2���k����t���8��+�F�g��UtL��Z� #"_.,����$�]�n��8�q�Ď���k���]��	��o�b�'���8޾U��efg��l|nt;����Ք ��Rm�_��J+�K� h�T�5X��h��&W�k��L��[�J����D��+�A��O��A���Nϵ4"�I~���	:BX�INr��TX��ySl;�3q|z.��vŢ~.ܪ3u
(j���]cX��M0�W���k}�	`|�?#�&E�	��)wظ5�c$��D��^���GKӍ��#&���f�v�A)ް���]�oF:�a ��'�_�Wm b$�`��]*���%�+8��*�Ra�fR�*�+c�k�A�m_-,�L�Ա���8�J��	�����?��uNG��'3kL��s�����&�� 3)�b�Lnn?ͳV�l��HTl ��I��I���)fr�\M'�gËY�K��P|I��d�|X��Ea�!�l�o��)p�Cv~p�k�c(�����hxA:	����?ֲ;���YUK�VZ��1:���N#ED�P�!�x�\����*~��̲@�)�Q��0�uT#��G1�q���.�s�@�R�X4w�#��A���E����=�kF�����g	�"M�����+������E[����xx��/x6	Z�D������dIkr���Y�Yt�{���E�Kh�M�C/Bݹo��G����o�� �d&J���(���`�j'q	�0g�y%ۯ*#��vf���m�&Gf;0�;7<e�+]P�����(��ޞ{m�N��_��6�i����M3��;1\ ��Yi
2Ji��^��\q��Ϸ��2npAF�C�I���or��5sas�߃�
���}gQ�|&�Q�T��0XSltg�>y[�w0	{�6'��V0�9��h)K^��?��0.8a��+�e=;o��@\n9��D=��H����,���:#�4T�`.�<��ü���1��n	 ���6�W��;ȁ�	\�:b�~'M9{�� q� ���J���|�W��T<����M�Ñ��C�z���bcG����īZ�/�1?Ω�m"�g�Rv����9qg)-`�y�o�1�0��Kw�|nNh�4��'��;8�J.o%Wc��pl����da����fK��t���jX�P�H	<�:L�ml��aH��B?��.��+����^���4�ԍϨ�[�\�x�<���Z�&Ҳq�(�dWZ�j��P���	�Pgk��-SZ"%�lܑ~w�Lt?��L�J�'DG�]Y�Q�󧚩Hi�LH�:@��������ص�Y�w�nς�X�.�ĝ4����i4<؁29t�Jr��|n� =b����6���qD,?�{�IM>��υ��S���!��~]����bJ7I�K}I<X�<�y����o����l��4�UbL�!�its�:����U�NXO���І���!��W��+��%��F80LL�o��ql�+�É�2Ĝ��xI6=��"�KCph��Xr�H5ʍ"Q�b�Gx`F)�^[k��*F��+��`&A���
�yh%.�F����T T��n7�ϣp��p?���zދH�/��V�f�J%�I�!����V.�0(�8pko�U�����kPzx*[/���8���`��\��`c���7�j 0�4C�%@�g$rU}�yfMk1���xMS��
/�$3.�Ξ�uP�5;�I��e�ԫ]��Wf�Pu�YT0T	2,7K�]}����P]9�K���&]�`6�Uw�k��J��^oy��r�gO�4[RgF�w��Ƕ�IK�V8���	��E�K��+tax���=�OC�6:0O������"��+�$�cD��{�9�xGXغꈹX����U��Sd�>{������s�J-n�F��aF�oQY�w%���U���%/��1Y��p������k��X�� �Ԉ���	k�~Qww�=����d(��eW�L�0i?��!ߚ�@�@??�n���U���֪<�6�͊��$Q���a"��Z�F�0�B��Y�<�Γ� $�n?S<DR���s�'���O� ����c���'tv�;��� ��G�+�-���n ���%�q��Y�2��pʂ�i�_��>uA���S����ɿ{����Ƃ,��PK`��;4������iK�d�Y�glzQ�ʊm�N��`$_����?�H~��4EcF ���>���)-ȧ���mpBi���!a��mR �J��� �l��ϣ;ʺ�����w~a�e'E�p��Q=��0?%�J������w¼@���4o(s*��)��AIX��o�pOc@�>-��U\�c	!�^��ת�/Ϧw�>�iY��Κ7�lΈ�R1Or^�!C`S8���_��p�Sς���j��B�)�tѻ8���V�y�?�%k�H��Uҗ.�E��`��R��d�IO��O����3�\t�_��WSC�GٓN��c!/���L�����fncC�q���h���|p����� '�pySe�������Q؂�s�v2�G���y�)�H8q��bЖ��E.�d���s�ҟ=�Fs��j�<G���A,�\ȿV.6Ɵ@������~�rG,���r9�D4������ƶ�3u�Y��ځr�A�	g����9��E�,�ҍ��r:�:q;�Cxr�'(Rn}埀{��8�n�$%��5R��xs�?�^3�up�F˛k��u0�/��r�&	JJ#�}$=)��(o�h�r������ۛG��h�U�5kH�<s��j����3��2O�c��.Bt*Y�J�\è�k���E>R��v��ѕP�99�.+���2b����o�HL+!��8}񈈌(.�%�Q�|���\d�ձ���U4X���Uqׅ1ӐG�ED[������M)R��A�[�LS���k�j�BK�������ؗ�t=�c+�M��C�Y}1�XW ���mϪ�Q���Y�ϣ=^C�$A��F�����Ρ�𛾡�(����p�gx�|�D��������J<�%(h�N���,�&���u b��9:h��䜥`h���Sʠ�#-|8:�	���2��uF�Kw��+	E���D�$.=�� >/z�G�u����e���6x;c73y0�`�1]EW6�{p�9/@2�i9b�R�]�L�&ݽ�2͇����!)�]���쭥��&Q�t��x�}�{���`F�lZ�J��ũ����)t1������<�­I>nt����3?�8&R����z3��Q���)<,~x#��i��f1�<���jI�I���[�5̓M�|2G��AӀ8��`��?� uV��庥��p�5�	ke��'��� "�>��:�[��	��2���L�#!@�nZ��j��)
��+9x��tꦀ8\��dO�@��Wp@}
;=۲�n�*e���A
X|z��;��er:o�юa�A���9A"�x){���I���K�$���NW�4 8T����2��*��dD��ފ�d_6$]����$>��Yܧ�f��{D�(�J�N}7P,��y�@Nj������*�ч<�{9�
��0:�!'UA�`z`
�i@�3Rݖ\���x��̦�`6�3R�7=�����إ�� N��g����L�z��S�h,~�LϹ{��8�8u�*���w���qQ��E@j��N���R��pE��c�b�
��k��õ�I�~y�p�̵����h�d:)��4����A��bD��3�f��뼟��_u7^I�D��� kEB#�)L��&&�<�h�S�2��K+֩�r�
ɤ�6��ޖ�����|)��EME�Bb��`Ʉ�{k�)�ڳ[�	���HS���Ν��*ky&l%N�/�n���=�� �Pf~�x�O���[�� /��B����||�&{��$���U���4@�b�=�����@%���5�!܀��e3[�h�駋�������_e��܆�
x!���k�#V��0�C��H��I��4����mX��:�{�O���	�D՘���k(��2�g�R�C��W��=C�b�?�&<t凤�`g�PmQ?j\��+=���O�a4��b�+�,6I�#�/N�'�;�WX��K0���2���p�@
����?j��"ZGZ"^���s�U�(���o���E=��k{?z*xXu����f�;D(�v/H?f���Q����=gU_��x� �h�G������c�Uj��y�z�;��B��E�_�@jtk��I��W���=/�5 BwB�6��]5S�^�W�6�׽���5bݦ &Su�sj#�JQ��T%rd�HP��	C��_?S�o��oˊՎ��>��LIo�}���r�@z��[��%�{�����lea|c���'��^2f<�e+������=�ͬ:'P��W� ��C\t�d��߂A�zU�t��mM�o�@�W�0� ��](ӑ�
>��2:��2�j��K.� ��t�x6�ڀ�{�?��i*	�Z�O�b<�֧bs�>��B8D䋸��63GX�%Fi�4[�3����$����ܞ�qC�ԱLD����vmoR�U��k�|u�cD	����r~4����^	��8+ř�(��_����4�j�*����v}iv�`��#=���Gw
t<���s�C�Qd��)����}:*E��C���H���).�T�x��� VMM��Э��z������Ņ��A�|�F���2r�jŦq�\�V�N7�iq�EP
�>��S���/��^
�){-$y(���ƭ�A@��h�}�3<p�#�0�>>��+p�u?fY�'�X>�ߠ���7�_���4���/�KU� y�q�������f�W�E|�|��!�`�t5�/d�j�'��{������a�$$���Ne�h-h�<���.�42E:�`%&r0y��5����1(�	4��}�C�."��;s��$�>3���]��Ib�4���4��8W���'�,��w��8n[��]��;r !/�)I�>��x��� �7x����b�C?��n�z�D�F�'�E��]q�g4џ�\�*q��A���aG�ʌ�Hl�bt�V�t�`R���@B!#�q�1����,3/L�uCE�VQI��6����i���7�I�D����' ���3�Yv9���7��\�+�9��rV=�b�����}����x?BI�8��m��G����#�.��	�gړ&,��_(�1���)J���T2>�b��Kܷ�S y��^|��m
7���v��c��.��5Z��-Q�W�7$�q3.H�����p�dCK=C�p�t<�wE��d�>0f�����8�;�R5�O�e#�$h�����
��tφƛ�|Ku
���n?
�
*�|�G�j:�ؖL5��yP\�l�2�X��^���wJ^C����G��pg�����xQ"7dyZ������؇��廬��������ep�O�NeQ��MޢDM�)L����4T��3ȇ�V�� ���K���`<n�2�,HE�T����v�!Z7²�5��MG�H����H[e�O�۵ς(ϯ�