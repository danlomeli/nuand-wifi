��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����xLM�����`,5?p�"���N��}߳�^'��v�Y|'�XR��f����mM�x�p�xV#ڇ��76{��)����L���h�:��+A���9ߨ-� rā�SZ )����C.��&0C]�-��[�3�-���+��պݣ�k�J�vo`�A�����f����u�X���v�=�а���]Q�Wۿ�߸�=_Q�X����j>��Zw�K��SvX��ƥ.���#�����Z�0���#7{��\S$��@1I�QX~TQ�E��db����۰� ���>0�%�9�j汈��}��1� ��2���h�G��SeY�a���	'<x�p��k�H`�H�j^y�0�s�78+���ֳ�`�R3dW��_��{p[�?$�s0��#�zS�_��bH
�c�p�IL7]� |����Q�� ��Rr���=��E즕2%�����`�^��l�q-�]�p��jf��Ӽ-f%H���ȳ�>��+���M�71��4_�) 3�46h�rb�J�W� k�h~K0�>P$�_n)���5�r�j��W�J&޴o��$>��6��ŀ�;A~<6P��K�~��f��*I
�Z��}`q���ApC��n���g���3��-�іrO�mF���,�$��@�BI�q�}��Ȥ֐����î�䂧��@������U���vU������ �T#K@f�㯁����|95<@���+�-�)�����K���FI�k���*@�m&���
���ma1[�2�u�I�\�U�yu���o�|��2����;�W�W�}P�K>%5�'�8���׫=����k��,�t�M�0�8]q3���N���GvZ�i�+ C�e
��Ќ�S�v<%���q��e_��
�k�夞��>ZO7E~��5k�TW Aod��eE���G���ɑ-'���?�G$����ќ����8ɸ+ 5ʗ���l�d��,�J�
�^�3b,�����J����#n�zK����z�&��;|�\�^���'e�W�����">�w*	FO�Δ��v�ƺ����U4A7�y�������\IҾP:S��ZC����8��d;#E���)�#8��a�K�C��=2OM�D�@`�f��J�F���Xz���#E�U̼���G� ��~N���ւ��K[}E�xN��x"շ��{
0-��5�5Z��!��>d�!��5�R�n�����nEV�@�����7pRG�6>0��ҟz��蝝���j��A�<�~j�L��)ֶ�Z�(p����\��5��︳����;D����NnMC`�(����\F=Cƽ�)����=FA��hp�=���]�2�OТ!�ҼݳIt3N����@�]|�z(��A�}�_I��f�A�a,��{���ˮ,g`�-��u�Y��r<�y?7Xo<L��~+�Ѡ�I��"}W��,0;���{6�@�<IF�=Y�"{R�ҏ #���u�d�ɞ�O�L�A�&��va�we`2��r�w���-�kq��%���[�ɳ��KK�'&Y��a��� i]�
d�O����OZ#ZP���׽h!�\�_�Z�42Z�VB����F:�&��02`���<0����;Ү��reW����6Y�DC	6�ȟ*��i1���	�Ͷ���(�=�9��[�3���~RyQ����$N[�;s�ʫ�����_�u]�.�Q�"�W�ՙ��,��|�&��#���m��"��v��DD�{�(�;��m�V�k,^���w�GM��꿫=�B����"�Pm�w�Ô�rm0���Y�#v�^[�a�ea�V���u��n�s����3)ڒ>��o��p�B��4���1�\�8�O�K�*y�`��l��a�p�n|��ȯ��Rhg�I�:����6&;��i�)g����v�J��
��J��p�Q���$�_�4�+�y��qD��p!?{��3��������@���)'��gK-���ގi�r:\W�q���m�������B����H��$��x�3�����k���T��C��0	ŘV��L%�2��c��&�)k�]q��׵D�ޞ[�/���18�{���
#���=0�+h�O?�5��G�WQ����6�bM��.��o_'�*H���{s������$�<�R�+�~(�������o_M[�`���;��s΍��;��U��0%�Z�/y�X�e��8�!`�csS����U7�R�)�m������QR3��#�cV���riKeӧ�լ`���羀��
�D��_.8�q���O��ʍ�^�.؛�m������F�wr�^��:��p�T�9x�hK�p�>0\�^ݹ�(<�a���Pr�{��tE	��^��AxQ�S�&8�db�8i�< e�,/������a�$��&�� �qz�Ơ&�L�v�)�!ld/�[û����� �䧄@[Qf��F��C���;�7d�C���?JP�����������@��^��	?O�p�Aޔ�W
~V�W�4��N����H��ex�}��q{��	7<C�4>|����6� �9(�VT���Ǵ����д���P�/�d}>(��Hב�k�f�Î���,il�C�Kӗ�GvK ҡcK��j����%��5��Gq΅R&u^���1�^���O B.��&x4Hqn�8t���0���/f����t�A�<���N[�ڷ1Ϯv��n��b��}�n�u,�� ?��_�O�����	V���B
�?���;�@���s����?Lᦘ�w�ou'���ۦ1yGM�ϝ��+#|J؅��+�eJ�$�_eD��d:pfs�����jl$�V8�
�ǃbV�1�����d�$�;{-^��P�AER������*��I?����щ$e
z��E�9,�]f���%�v$���dh�+_.�>k\S�v�F��jn��h�f@L���!��hC�;'�;@uk�B�Y�f��&�Y
K��u�t�՞\���J�dB����'�<�#�t��j��-@G9�2F��j�ߺ�
3~˂����GM�QX�|���������7[�^����Ao(�[��	C=,@�1NCe��WO5:~��t���
c��O����㼳�>��y�nP�j��Ѳ(��AyZ�Ϝ��i1��fu���1�ꠛ�/�XB�Ue�ك�d3F�E��ƻ��e���@���=@�)�
V���{;��!����r��'	��4�&�&��MW�J�D���T�`5ʬ=��k��J���1�Co�I[
[��:�k�.�����8���|���\'6c�M������ .�6>5�C�i�0��4S��2����@��F�:�͉3b0t<�c�8>�Y�=rS}�z�=R��Q�. �]�8p�P�Wܻc����wN� �<��G}�X���Á��țZor�Y˛�!�&�gY�T�#�?�W0�m�B^�X{�U����%�8�oӧ���tاJF�t����F[�|��2�a�ʽT&}vvX�N[xP��+l�
߄�@O�x�䍹o��-��K��d��#]kMIE�2 ӫgr=���
�П�=R����Hm�,�wɾ�0�� F������oD��N_�Z|�^'*��� p��H���Z?;-�����Rp(���=;*��n�ې�%ݳ��7���F5�����?���Ҧ�x���Þ�q�+ԯ�߶k:���?���2ר˭5��7��������f�!�0%�~*�����XB1	#r�ÈM�i��[�erh�u���e�o�ڰ��}O���^���\S�jc�#���^��
�:�c������,�*�v-L:���Z���\_��_��,0�+���,���v@�^�l)h5w���uL	��.��T#ty��o��N+�;����*�ٿ[�P�_pm)���Oh����4cg�"%�Z�i@uS�١�_��mQJ:�}�^c�U��B��$�]e+�,��=�G��7+M�e�,��ȴ�kv�ȼp�h�%A!������r�Bt���;E:9^��;N��.���z*�г��df��E��s>��pȢl��(p�A��.�m��] �́����(�?�;P2�%L��i�3�l��z.�
��ŮM����XlF7dZ�ױ��M$He}JX� !cMKï�7ݜøֈP}]ŝ�~��\ x�H��6Kϼ$Ӕ���<ԯW��_PKJK�$�ch��R��v�
�+��sL�-6�7�~��׶Yƥ�@��Ǖ�<2��1��E7�V����Hk��eF��=x�"df�e��K�s�������:�ߘ�M�˜����n)�%����^K��@n)����u��L'��.�Q5�V�;�,;M���'-�۪�7�z������ݪҰH>�s:o��F������
�V�;��0��v+����-T*�B���im2w�AL�{?/.I�ќ��d��I���~G~Wߒ��.���5�̭�*��P�y���J"JWWE1�	�ۃT+�f1;�V�����#?��ax�89B���a�6���	�1Ѡ�6b��2h��Ӷ��ȉ���V9�d�xG�1�W�#y�\��g=�ӿ{���\_�*���%Q*�?�����o�ǰEdK�ڨ�f������l�7h�NN�9�%N���J�q��q�e(/�G ��[[�Bˏ�c�<��T��I��ӗxjq< D!�u�P질+R���%��v��2b�c�89��kI�j�>����$Fa�g��t��Τ\�@2�l\xR�(?�0G�0�S�[<�Ĺ.g��4���/��{&.�k=(� ���E�͊�*���}w�;�t8�XX ^-�A��
�d���_b�[��R
��Z��M�M'�#RV�i�+G��.t�9.��y	����[��_>L/+".S��Ư_O��̆��ߊ]MRF�9��}�	��~�e�6߉�O���P@=p��ѯ�1���i���%��G�p源_�xW<U��=��!��M�{���)`�.�S�c+[]}W� �/��z��������]\�4��)Nڙ���������$ʏ�?��S�pjH*������a([18�50 ����2�<O���G�*���{L����f\	�)dx"����xnjQR��i�u�X�P�_��2Jy��ˇ�ٳ��1j�'��FZyGxq2�$+�6$�����-�Z���S���8EyM�nt�)C���Z���I�K���.7�*��J���☙�_3���$=*�$X���B?_7��I��0F|9g?�mv�7�1{�f�jǳcX�b��F Kq��"���[�?��%6�b%

$4�h����?���G���K]���I�b~�@���M日����9��Lf���}G%��'Ѕ�v'5C(�O�]��2^}]A���.�Ѭ�Ю#���-W�ժ?0�Y�� U.Cx+��!=rf?rZۡ�����zE��]ACĨ����q߹�xJ�CE����1�w�w����b{0Q��}���n5F�ɯ*�X�����-�$,����ª'��Ҍ���ste��A��F:�X	�UQ�D���od6���E�ު��|B�a�B���2z�tۗ�{����^sULuv���^��(:�szJ�6�.k��h���n"�+��.5�,cB�����ȣ�;�I�I����!S	�"AIKl��l��nKВ�,�I�+��:�}�O�f\�b�'!��̫I ^�q�Q�G{��ӟ\9lK�s�M�⎻ϖ)���5Ŵ��iX�1�"c��j� �_�[���V��Wr4�2�ʱ�.��񤡛�C(����Pb��G��H�u �I&"(�e�����'�{��|Dc��b��=���߰�k&k���q:����.l?ե����o��@&���~b�!��b������N%P�O*�*b����ۯ�q�m��*$����)o�Eq�6���n�	�����,Nw� �Z\�
�H�Vv��&gTzf�[���3?�J�"��Z���4�Wy�._E)OYX����7 amx�C!�S}�����M����O��2w��p�*L���U(V�~In�ߩ~]�5"��b�Z������x�R��2P�����L�`� ߇(�o�;���t�,ݹԑC�9U�gH����s�pT�s��MC�c\}=��E�J�`��_-�'�Õ�f�&�jO>�B)�CyQ�Ջ���� ���$�w+ܛ�u���d^�v�D�
�i�]��Gi	|O��0s��pB#�A����ޚ}<�i�H�������<e47gϖ&"`�r��G�R�5OsT�H-��W��#ԟ�?���`��lV0�(-B�R����=�0��ox7ћ9��HSU��2+��R�k�y!�{[L��9X	F�)��q�h��]r^��8��`|�uN�~�X�$瑷�).��:�ޘ�9�8��c�Ů��{W����?���Z-����@�-��kA�t���gA�nS@�}�۪"?C����[YRK+�����.�6�?��k�
r�W`S��q��ry�Ū�lw��c3mX�4�a%i��"�8�hf5��`jt��y���ח(1Z���Ln0��y�cf���"]*n���P(�D@1�����\I�F���x�~�8ͶLѬ�Ƣcx�2��_*�ê����z��x����#�G�1�S����i��+��dOSBk�p�)]q���x`�o��w���>I��y�򹺴9ڿ�׃Ω�J�z?nt5a4c|j���� ��N�9��`�yUTF�2�.Yj�钫��2�D`���2�o��+�΅:�Jf�f|w�D�«�:���4�<ѫ�b���8J�ٝG��q*MR�e���I�X^��G�]�uʭ֣����!�χ�dW�^5&w�w;��4���R� �_6�ċ'�h~QC�!E���z��_Պ�h�XN�{4�A�M�I��)������Hz�G�$g�֗�*Su�)P>4#i&���5)A�Y��3L���m�[S��@i�a���K4�Q��W�/dhz��ՠL���
��k��E� 2K���`�2K#L3��E�p�+��w�0?��L�6	� �=�-	.58��X��e���;^���LBMc����hIN&��&਀澠��N�­�Iu�?u�)'���?�%�Pfǔ�S�!f�*GLj=d�F6^�<��`���㧂�Cib�����Z�&VU#�����Tԉi��j��(��-�[�����9��:������X��/�\@�h7����l�����K����V���{l�0���&a��W�%�J��8�*��l6��zrw�Np{WY�h��#8��ڐ@SW�B!&�p�װ��;M�����Vo��iX�� ��bIC`����gH��I�u��J�?�!� �f��}���J^�J9�<%�����>\�I�i;���`C����ݛ�3�C-�����|��f@G	ν?�����73f�"mh�py�>��C������7�W�'��;��s����9bE�'�S�{�n������K H��8�Ԏ�<��(�&=�H�e��/�$#��@�#�|��ۖ���Sq����<5��N��S��d-�GS��9�/pZ��r���:��3��8{�st�e2e�}q�����K���h��K�Lx�Ȟ����5��㺎�C.iv�\�v�N���X�X�0�����*��+*�E!�F�W�O[������>�ݍe(@h�l���x�q�4���W`8��zj��k>L��'2�������M'YP@r�	<���,�f�W������3�>�����n�^�Z�I$�T�'���P;��/
qbPJT���_���>�,�ve��j�2�4h�ʜ��aˋgY�`�J�Xn�����\��fZ��O�M�1��ݙ'�߮��-<J�a����t���9ygfgY��3tS�vι�VK̖o��o7��Ԫ5�[���-~��*�v{��(��W!����X⸻*^K��u�?BXb���k#����[�S7���\��}���Pﰦ�2ǉ� ���/+@I���<��N��n?J�_y;����ڦ1x�n-��;��}��r�=9�?[����i���/3���+�)IU0�\6�z�S	�ޯ��ɸB�K`�t���yiٵ��%��3v���*����lIy���.���utVH&xP;�FE�xG�,|����t#dr�����p�����0D��{Lu�2�Za��a���y�T\�� $���4~>Ğ�W���Ҁ{���C�y\��[�:�1�%��e��3��t�&�B�~�Yu��Z�4RL� Y�G�kv0�YDb?��B%[�\�XR]R��ǧ��8F�ER)׸N&������nq��v����q3��3Dj��!��ɘ�&�m�Ý�N��BU��+�������'Qr@����;t�I�a�|:@�����AU��zSxwn��9�5R�m�a'�Ѕp�GlO��t�̎��JX�� 5~S��� ې��m�V��r��&�2K�1�[#ң�R���5^�W��~�X��YD��6=�Q՟
�a��اpѡ,X�7Pe��ߛ��u��C[�}�.���?�meȢ�B/~Ji��_�Eе%/������mPr�����NC������P�?f�K��n�������Lڐ&��(��'_�)�ϏX�W��x21��s=F��`�P�[e�@�_�g��&�q�䏒��
CwI�%�]�1��'���r(�)u�>nh�E?xI�\K�:%��
Cc�Nﴚ�H�2T�{ƒ��01h�:�����Ϥ��<|m����?A�ֆ��,S��(������/�k���Q��5>��_7��a֘[{�Z�V���b��(�l(��" 4�g�|�;m �x2�+�-<�F�͍V+)���3c����p%�![�(�kF*:��
N�<Һ4"G��/�-U�a��3�4�ĝYԞ�<������(M�IZZ@�~A�
��2�sy�߾���U��G�E���bT\�JN&C�\�N,)����>��A�/TS�ϕ��;x�8������5��M��!��f�lB|"��VTv%L�Xk���/��_dBch��dr
p��'[?�a��YnBH�ˀ�R�������U�C��UӉ�+݉>�жfT1���T���f|�Mn��J��	�*@�����S���+8���:Fu[����2���:#l��`y��niN�e?��>il℉r��f����T��/���&��{�E��|�c��^�?tk?]�`*ݥ-ܺf��@��Y��9!#!�Tےo-�}�l{��( �QrR��oJ3�v���CP`�����P!����O[�dW�3tx��8���x���6/���@ֻqBh�����`ղRq�D������ъ�x(�,�:��� �I���Q1���+�|b�+���}�2��V%{Fp�%Y��%��|��q���x���[ �hm�k�����P�)�0Ly���3O5s�x�L��h���s�zg�����l�Y��D^�s�"M��6�ߧ� u��eR��|U�W�|㞈�5��;n����
?� F���. CU��Rm5L�����bI�9"s�eF�' ��Μ�Y��0i����'�d�KK�Ң�^̗s8��&�,>�[$*���� m���?������Tl�T�q�Z|�N�����տ���T��ۓ���Q1��(��)���VZ�	sn�'(Z�z��e��W��o�=5bȺ��<�4f���DFH�s����G��Z��ݱ�� ��}��O߱e��YC՚�m��d��k�UY�C�'����H��է8�o���ᴏi62�{�O7�B;6ʻ �|��yD*Lx�'M�E���j��jX̝{��|�Dl!
����}�%<���+���G鍣9�Y<��6�< ?,�A� G�,��ab���B��"�|v��d�`�?*����B���X-T��ZM|����z�y9}�LR��T{i�)@�T�D�씅��M�		�q��w�� �p��N�wc��/tw��e>+�9O�qEr�|m�<�����Lꂥ��K���׶�]��fyb�_F�el@	�R|:e��T��q���h��J��'T�Ӄ�&�)��ӈs;��L�Q#��Ȁ�s�"~�Q����\x�?-��J�誣:�YI�z�i��k��5�E!� NAJ�<J��q�M/|��c��9�DV����|f(8��i���ؑ��-D�9ˌ=�����^Cϒ�Y�|�T�Et�����ڍ-e$	.~�P���Z���^��l6��ր^֒:�兔�ѽP�;��u�*�R�Q���{����Uô���X���
=ޕ��ֶ�9�$-J
�\�n���՜oi���D�hA@N��ʨ�ʯB\�0���E����P\'bD͞@�%ئ	��	�;?mBR1��6ǥ��K�Y�}l��؞���tj���<먿��Ja3]��~S<�ۄP>�� �'�H���B�ػ��e���l��	ݓ���wg���V}=�A�V�B}�^0�3��z�bB�]y(F����� ��TD-�9����Q(�@������!0FS\�tT�q�c�O�?2�h��"ۓ��6��4;���KH"�ͧKle�b��dY#��]�Zz9@�/H�&�M���]�rnY6��0=�	6���O$�������'�{+�k�����~����\p�ƙ\Y�e�"��N���� �!����p��Ř���^@|�D�y9�NJ8y��(ا���
VP���	{$�Zge�����EeE]S�%�Ʊ(�����6�: ��x���m2ƻ��]�%�ڋ��+�h�F�-����Ƶ�ln0 TF�"���d�q7ASM��=3�hV@Y���Ӌ-2NȠX���:2���`��OB,�q���}�3�B�}4K��f��5����*��+�%� Ꮵ�17���f���;�6r��X����5�e�2�x~]��Prl]Q7mG�2$���"�]3�Ҷ�+�j�8ޒA�p���տ�w��c��m���Fk7�sb��K�ڲ.���T�gD��A�Mf��J�^�����%:!��S����q$3ʧ&���� ��L���	f|���rM��Et���T��-h�V��sТ^�4��n����ffN�m^;K��np���R�o��/~��t�_��} ��A$@cKmΟk:�]������Q�������X��du���
��K�ſ4�,聉CT+�3�״0k3�D�O:�)t�M �L�*���S��˄�+�ŵ���xM�h�z P��ZR�*�MQ��`Q���{�jhl�GSɒ_�<��DW�3������ۄ[��ư�7�ӝ�~c�*.=�R���Q�'�Z&�S:��v��|ĒŇ���WȰl�)$VK>�� ���)n�+�\'�U����$>��q�^�|oX$��rq#Rl+���Q��4u�%h��x���xǞ������=v۴���b��a�)_�IӥIoI�"1����)�.���c��P{�gW��EpNY�*�}󚯏��j�_��&��4a�ȯ�py��d{���?;�h(~�MyW?�Ӆ'�I��������֛&�V�#.�ak���Oz�/�.�Fiݨ� 7��������<k�)�j����{*�����ks��ԣ����;�O�a��nnLm �w~��g{��>Ř#4qF<��q��]O�2�u.8�UB�>���-�,1 ��C^�}���C��P*���s�L;7t�z�p6�j��	�y�6�3B��?���D��/���b+�'d��c�E7���x�q	�gNrS��I��,�_�l7�	te��e�B/���t,7�rBR\�L�����G���D���{x����Ҙ}qq[����4c���!��m��,h�� ���@��"��!̉U
��t�%ET#� 3;�$����PC�'P}���S��h1T�Ԣ8׶�g���[�O|�������l��`Lj�T�^/Įckn�Q�I�(��9u�J��H��Jn�P�r�O��9�i��C�f�]̤A�
������!9��LI
���+ɘ��7>1�x��B��J�2��7�Co{�d�u�z�Tu�4�P�Â|6	�?�i�;cG&J�����g�xm�����|�q�b��<�n�:G��	�Jⱡ�.�H����0)�a��J��⮂��V���?<��WAh���K����L?_N W�Q�kN,���ã�d���	�m�չ	�
3_)�HY�H�ֿ
���	'�����7�g\6~15�c
� �ö���š{����$��Q�-�����0�$�Z�Tb�GT(�s����]�x3�:j�	�W�����ĕw`}�u՞�L��֟�TXxR��},.762Uӑ3���/�Lq�����7�[�S[^ �-�Cm���E>���n��s��:�5-T���"��Rf��ń�5�m/%!���ɕ�M�<�0����Dk���M8�z��K[���Lf ����\��9���<����TAb��_҇�?��b'��S)ǉ���`��{����4����s�~�'�6x5n���B� ��v,ǭ���}$G~;.Z�h����Q뽈F~O��*q9��ϧ�;��D��/v# ��p�$֎��t�dĎ�[��F��q����l��xk:s���C�\d����pc���}�}:̄1~�3���7HW�](����!>����()w�}t�þ�7��/�LZM ���)��v̒��RX�T�2�ǚ�?A��P�
�������$p½���X��� ���ҷ @�N' u�F�ԕ��61��('��
��Or:�"�s,I�?:k],��]\�ι�Q���WR�Y}��qm��'V��Mo�����uh��J<���bZ��ԇ���BZp����U�2��։.'��1�V�V&3��8?z��Serpx����m����!FW�/�A�0	���MB�ŝU�k�语>��`��Ea�����j��K�%�	�:`��f�cQ���S���`�d��ч��X�E=ׁ�(J�ˠ�s�(&�\�
��a����r�A y֮2��tjnͿN���0<���T�_S�!�����7�!o�qjݣ�,��Q�c�߼��q�r����ŏm�0�l�Q?{>yc���4$?��w�X�^��$c*o���n]�K���<G�:����h�M�����f�TO��S���7Ш;h��FO�%Ӓ�{L�\�!9p֔ȁ1�[~8�+G���R�qh����3��x�j��J��!i
�2�s{P�#*P��7����OB�Q2G��!�;����;!	'����cXeC��Rpo3�4��Ë(p�l�'�N���y�����m���B��bXuxf	Ŕ~\W�X�C���anS���pV�9�}�r��o���_��!P��I���m���q�k�h�	�=�#ѝ&�p�^�k��.��"������_�]��!~q��O�uw#��^�������	�lg���C��iRSL^�O#5����	�8���Gh��Yu��@'͖��42�P�T��ߗ�W��A������jzDs�q�~��{'w���;��������f�n��2��Rd!���ߓ���z�Uׄ�b��6� <�����ͲK�ɠ*b%6�z�P��<�#�hs� �6x�����Ƣ���ad�ÑaL�p�'�����j,��|˹>�jJ������&� a���3y3�������[�d�o�U�P��X~����������i<��%�^���`{.]'�d���s�KQ��f�u
%������oG)���6'f�O�l9u��7�ͪ�Nܵ�!��Q��!<K܈	��[�]KC)%o���#l��	�AI�������KN��\�k�M��Bz��#�'�Ǭ��e0dC盵�v-�����:�6��~��m�p�m��D1�'�ԩ��,�!�k���qcD���\�6��z���N��n�lȞ6Dl�ze%gDe��su��G��j��r��M���&���z��e�P�`V�>�T#���oIM��i��KG��<"5�1`?��R���!3�����s"���`�;�Mcw�i��`�Erh�`�{,�)�b��V�����'_�
���G��ز虻����L�5Y�>��c0����QA�Q�L�o�TP���Lcʶ_�|�W� �~�gԛjE��{&��\��U�u�bx�U�6��G�b?�X�h����7FZ���Q����N,�v�T?JN]7��{��~����6���' �dXyV}�t���q�S�gv	�[kn1�=�5̎'�
�n)��ӳ�C�q��ţ����.Pk^f�o�K]�� i9��r]=K�$�ZT��sr�P��@�q��/Ry�w7�Ź���r���i'f��]��iJ5m�{�j�1�F$�긤��\n!}9���gcփ��=!���<m�b	�飗j����{�G���*}�Le��s�y���H3�V�����Mp?��/��/+�=i�Lc�qe�sQ�TY�m���{��DG(�n�� ai����h�	y�H5�v��-�s<�T�]���G:{XTF>&ȫyUT^�?���޶�?<��ria�;����뿑ڞX)��Q�#��X:���M���HU����Ǻ��2",Z'�#�K���
��~�����:ݗ3ٟ���Bj��o`X�}o���Ʉ��A�GI�c��>���Jkሻ�d�ug���γEI��4�ߗ��d1��@T3&���<�tl�1��z�TS�� h=�03CA��|���iw�EQ��q�1�����fO�� ���a����C�ϕoR���i
6"oYc�a��Q|����ԝ���Å�]u���\/yl>��âAd�I�N9����a8#���`��:��~.y�����Xz�>���a���P����w�;����D�����R�Hk8� ���_{#�=^	W�Cj&L�[;����Y ɜ�;f��i����L��m�>�[
�d��${����݆�^�9�����=�!@?�0�	��������LIL�s/�P�a=EA{��b����w�;C��PB�+H"O,���Ó�B>Ha§�#����4D���� M���֞�~|��[�|,f7�R\�*�J���r�ۉ�X��nz��s1���j�~��ply�Gטѣ��M��̫����PĞ�A,��ċ���[τ������=�N��T�i�Zl��CGz�t��ǻ�_�D�`����R)�Y����h�
�b��L���V�P�	&�Xۚڏ9eS��e)�*е���>�F;��7�N&�K�*�ō��bU���{�wBH����"����_n�����h�߅RD0D�ka��p�~�X�s���g��d��1�k�W8��Q~uτ�W��m6A�W�ˣ�z�����bYrX'p�(�/�*]��uqf�愅=���
�ic����݀��`�hl0�}�қ�OW����+p�g $�@ҧ������E^*2�r�6aU֦���A�z�}���/���t�ʽ�M	t�����������pUSl�Zr��� ���U�@2f�ucX���Sߜ�i��	�B/�er	B�*p�%�C�L�_�B����i�T����S��ͥ�=�/�Z�ڴ�r$S��syXs~����1�㈒���|��껹���{zfi�bb��V?WN�m.E6��@�- �	�9c������F+�����yUi=	-"|� �$z(Iv>��� M&����),��s:3_�����WQ��Ŗ�	�)�l1<#�?I=��_��>��z~�_����/!Ug/W�s�U��}>]�M%v��y1�c�RD�C6'G�Ɣ� Q�$�9��t��d��T�-Vǭ��y�Kndi��ݑOKn�b�}!_|^/�j?OB����5xR{��	�3�����B��(���p [m�Y��$��g8�%yH���r	��ז�Y��:����Y�^wX�Q��l �@�׏b݈:THO��MJ�C�`t����}� �z8�Q��E�7�Q�O�>G�O�:U��q�{iӭfS%��*D�y�4�;1�hc�$�_�r���(z-_�;O_�.�K�BBCߒ��7���c"Jnd�t�&Y*��7�������9��}�r�8�F����^�W�o�/Tm�Cꔣ&$��R�蜣�Q��(�!@�W���`6��V6�O�Z=�2�]x)9Έ�*�5����+��*�k�);�|"iGw�.`_{w&�H+�`�+�aR'�g�b�ỡ�f����,�C�j����_p���q��v�� �X�",�W�h�P���gkr�uf �'�N��C�K���;�bU�3�V���O5]�B��������$/Y��ezT��
m�T�����5:��՚�s����'��Q�]ĕ���]�	X9 	�<&���4����7�o8�ڱZ�j��+F��g��~w[�۪���OUĮ+���ne+ơ&�B�H��4���w���]�
��5@��0ES`<�Ѝ�%��Q6T���i�������cbI#�J�S?�3�F�h���gő��v�MSb;}�$�ivl��7��{��������X���\�&�
��[���2���Ո��x��{����e�Qd~ʐ�:W��韱��6E k�z��uV���J�Ķ �2���瑦!���%z�Wg�)g��u�{�J?~R_gĒ~�:�!�h^C��S���l�LJ%.�W��d8ng���"��8�#�3��#�MK�06�x�����������G��L�������yrb��N5?&y�Fq9wv�F�qW�m{ _�t?���������;}��_n�Y7E��j�I�J�`䓀�X�|3��L��L�.���` 7�ߔrŻSz�c�����w%�6��+��vLM_������/��d����|�nI���A�`Vhw���{:V�=�hL�c�G4{���`���S�Dh.	�+P����l�	93.��N
�a�佩m�4�j� B3�h*�q��g0��6����f����fR���qB�g�7�pjA��^F�ּ�K�r�<R�b���ԅu��A��>n^ظ��I0�i�̏��)}?"mƳs<2���gT�2S���%;�6�<=4`02c�ǫx�K��~
�\���مk���s���%	�mL��Ј��PQ�)�LB���}{�OAM��0	I�
Y�1�b��%(Sw�c�t0��/��'9�Ǡ�����N7m}R5�qz�ⱇ�x|�<�G�>a-}�hg�?ְ4"T?Ca�Esm	j'�H�T����o���׫-�:hc�j^�-�ґ�gH�J����f{�H�/ |X�����fZП�u�/�=C�b`ym�MM=� ��nw)C���(s�Q�~�ހ����v�	��G�U,/����gP�锵��5�(�}
|������8oE-�a�f����'s�'�)�x�V�NnPL!ΚOX{G����PC�������!X�s-�$q6pP�XF�[��,�P*���M-�Ne�,�Y��(�2��z�#��N}�)L���~�E����&nz�G�3�涿�����*S݌�:�>��� ��i�!/���xX��I��h��$�L��_j��͕9Z�xτ�S���2�Ie!~�!���HC���Թ��n<���=��"�dk	�N��9Ӻ�����<v	��F]� ���V��C�͸8}t[+�ǐ*R����������j�A��{�e\�F%�Q�P��얎X����������X���!�. ��w��\�[1㟍3CD
kE�^����
b�E�{"u�,�<�W�.-M�a��
73c8�ۂu�����˽�&���@�s5z���nh ?��i(w��kwA+$�;�i�_��Ȏ��bkt�rLBeTr�@���U���jU�ndV0�t�R�(�"��{��.��JK�T���m��zX�z��� ��Ս���R��gQ[�¾�l��8*�=�����oV�B*����k���]�ų>5"s��
�e�8��[ac9����Xár��)�2f�U�����E�C�80�����j��υ�g�-����"k�n��J���!��r��5�'�5���+����K����B,�	�8���$S���ӊ�����uY�;�=Y,K�G�֪�'������\S��+����N�?1k�T|Ʀpv�EXd����r��dw��M��h����M
C�������$��������fYV^�57�]m�fs�fNn�p��nJ��z�ܚ��ÊƓ�~�����Vݖ����b9�N��\�2a�a�
u�d�0�ݴ��QJ���&��w"24m�����x���N�f�96��^TP���zT%����fI�jQ@����TκpTf����`us�.n�`�\�f���Й؂?�8��F����}sP�}7��6�v2,J���J���ʜU+��*}�z���)�i[��g�B�4��񑌅^  XOa� Nh�u&��#�����͡K��?� j��T�r�kC��1%���t�ŏ�5}j=�	Zⴈ���k`N��S�{�ּY{����c��N��Z��6���ii�,f	V�L�^| ��� ^����b�UK,��xʹ3����x��>�t�%؞Y��w�m�q�c��
ϳB̓�یx5����'�p���ԛL����AÌ��a-�i��F
�2�[�v�E��/1�!�}�����7�x�W�-D+(����Ng����Υ�(���es�Z�G�j��Q��%� )T����2-.AO�/J�]!��7Uvl(Z��h����o}s�FW����Q9�M�lA�E�'��T�k�����hd��<m�n�qK��YpԶ�C�F�D�KXF'�ʔ�*5�:<c�k��y�5р.<^�r��G��p���+�~a���|[�^l��9�Hc��W͉$3�E��E`�.*)Lc���L�4������x�_�;�l(���:�Z��(�X<�q���Œ$}/���J[~ͪ�9-�e#{��ݍ'F�]���ʫ. ���&j��l�&��J� ���9����1��"�� l���,�8�dΥN�%��	����At�dI�Z{7����"�^�0��Nn�O.t�%`�]&��v='���[�T�S@��I��f=7��`V��\�;M��j���:�ݔP&�\�̰��0���������I,1\����zf��Ԭ�����+B��M��]5��Y��E|L)D:�c���4�D�x��D�����F�^�!U��jBCqѬ�[¡�&�6����;S�1F2 Zא��B��EoIez�?�Tz���yy^Gߣ�D&QQ������,J��V������"�4����0yՁi�ZGM���^�C:�$ɌV��$�=�K��X'@"� ���`g ���/Rh�JQ�q�54��\み�d�[f:;k�z��S�˔ٷ!#{�]���^sLI��a(u��ҕ[��rre�I ��x=Z��p�Kԙ�5�7��K^��Pd�"����!G�,`��Zq����ޮ��Yf����珧^�T\�;��}�c�ú��S~X�_�L
!K�V�1�s��ioK<ɠ-�A%���tq(1��<�H�������n�hhB�dp�b�Ҙ<#�-=1�ݲ'��vü�ȓ?���WK�H�B����.�>�Q�oq�p�آ��d%Zک����n�_��Q�����7� �PC*o��Y�Z�ŉʹ�4�����t�(��Ih��yʳ����`����y7�[�3���y3�h_��bƋ]4CK=?�L��\<�2I�%zm�G(#O���T�T��t���r�T��m�JH�3�p�K�,A�V�ʩԍ{��9P�T�.�!­b�x�n����ޢ/Qkl�_��<K��ӓ4��`Hl;ll$�8H/���]�����ԅ��6р1sH�y����!ޙ���#H�)ߺ�)NRn����9p@)�������;F�˫$�7�<��Aҟ�8㖐E����M�	�2�����8P��F���aWk�G�qK3fN6�gX��GY%�@�:]ڞ(�	�Vuy��3��'3��ۑ%��!ǰ%�R,,�u1j��4nvO�6��
�H��=�<̀�|]+���{O��
3,0P�k< ��.��I&�9K� ���%�ܡH����/��ޢ���c.gr��Ӈ;3ş��q��2HH�4�X�bz��H6�_,`l�͜-��Q�x���G5�SC�5��BH�v��@��"��Oˣ��_W�8��ɓP`���<�H��$2ϙ\��w[f��xr�u͕Vz�~�Ҵ?`	,wl�'�j]�{͌�:��,��2����/����]��LN.�Iߞ��N��v)����3��}0r�p�	Q#?���4*]���Hx�e����w{��IH��[���QS��|�BحT�
-vL���3�I�5Ћ��ҿ�W�F�)�-gwrɿ����)���&���7⍢�g 2w/~��Fx���e�Cҹ�0(�Kyz����-݇0��`��/����n�ZסA�!<�9�ꨑ4��Qt����cb�Y�5���Rg���T<8��!i8�����w3�G���%�I���&�=1���������
a�����n�3�{���7�����(��z�Hϑ�G�of^���}�/�!�y�Α��"�)=��P��h��:��N]\]�O z���|����s|#FD�i��-�:u&'��lL� dvtf'�0��\�4F���w笌F�]�5�S�RN|'��L�I��$&qt~?��W5�������?�����uG���뛞3g;,���>���X^k�ʪ�!R�~�+{������5�h�~�A�������Pǭ�rEC
�86D��#�$�@X�E��e1%�i���6�#�X0�'�����9�j��f���ѵ�" �Vq��-����������8�]{LӡQ��JP8#��(�S�v d���^_�2��֤s��<��#��b\��=� � ��t#��(��Zj����7B�5&v�E��`���{���c�"��gL�7QFT}w�	���q*m�s1��×M����k*��Op|�d�#���l5<�6_���?����5�$0ΊIB�pa͟ޝ5�-WA+��u^�b{�<�<5����k���bl���]8�:���7�"=�v������j`��?4	�4��K�H��Ww�_'L+����pU�$�nI�"/b���7�����vڧM	�2,ҹ��ZHq�*��q@�"4����M+ ʹa�?N�X&j)�]�E��K�(�3�/�>挜�st�lڙک��&a��ңW6���Hw��^���e�D���{��!?�yP�~�s}�B�9���l�v(�u��f8z~���$G���"i-�y0F>���u�=�����D}�#Gܿf~k�����#L�Fa�6)��ԡ�(�啇��A2�W���˃Z5����t��'�盭�=2R
�"[�
���T$#�ʸL�g/�Y�]A+(��q�xwY��(�������ڹ"=�ʈ�\�� ����3r�q:Z�˫g�3� r�9sO��6�H�"��Nb�*v������zBBM��Uz�Nc$��^-�Lѷ�d�6)��3���O4���G�'�Z#�-�(��삀���Ϯ��uR�LA������� T|½�wL>k���%&�K]ur_�G=eCw�5r�m��$[�A�fV�"�~��@��p���U��d�� ���n��mlW~+�=:�D<�T!�@�����C|�~��ew,��ܳd/�#�?�17Va� �	�^��FQĄ�nL Ԏ)�X�L��J���#I����Q_�iϋ���-��x��k����&8�i"�b��n��Z��@�[+���"�ĮD�Ǟy��]F
����`�>{��}=Ą����P�1;��1JIA�yt�-q�݆/�E�*���4iNh�������U���چ�#v�����x�I���D㚇�1�DE�v����#�4�cv~|�-7Z�އ&�&
d�vT.�7#�2)gn�9+�~�B�^���X��zJ�E������W)KJIwBN#1� <����/ex��r���ؑy9*O����ꑰ�k�|��N'�tT�6#|67h:����^�ÚN&����sl�[q���<���ggZ�b���W�e�l�/_h3X�GS��p��3D8@�����u._��8D� �]�adpt ���IW> ��F)�W/gb�aǛ6�x	�e�sR�K�#�>@0kҸ_�1X]��g��ߥ�&s2� `�b�Gq|`U}�����a��@�b�j�q�Tb�Ej����r�a�������A=�3"�����-����Bn�S���k;��j�	|&)jS4@� ȋA�<�&��d�å�pP���,)�������w;Z�az�&�E9�kz�[�u@ ��Djv]���Y�˛J¥ )���K����rC
�g��A:�ѹ��@)�
�ۨ؟��&���#��Utu�E+�'AT��fb~a �:CNt��3bغ0Y�����Д���2���ּ#{�����z��l�:�]����nWl���UēP�}�	*5��ڜ����|��l$\�[��N�^"Kk3h��L!^�������#
B�� ���`Su��M��/�a���J�Mzx�M�K��Dv��,����|]U1��8mHV�S���F�_�1����ц�/���6IA�(o<2�Z�%b��w��)b�[��g�Չ�8HH��i����/���_�һ$I�+�G"�xZ��%Aa&K�a���k��!d-��b�R�j؟�e����q��_�KFɫ�AW�qKy	�/�].Ệ����ár���)��N2��ѿ��E����%��a��Y��H�"��i����nPԐ���}K�]���B@�6ͰH� eŖ;���ZW����Gb����ҳ�w������HpM�vi����f��*QBgό1Sc"��x�<Ȼhy鑸���?4�y��?ZCR3묈�0�P�$z�Л��f���<�$��a���>���0`
�Ju�^�b�>�
����Wڮ��)t�l���	�q��9��-ֽ"/+��A�. ����h�${�I�隟�������nQ�{6�U(����hi�s&oO��o?3�{y[�p�otoZ;����{��]���EN�>j$���uF��7�jΰ�����ĭx݆WH�2W։S�H�6�_6�J��z�wr�:�O�:�"�A.����V�xFb�oiRL��4<v:^vUߜ�PA�N�	��IѦ��j��$�AY�q�&������e[:�lحyfD�����ȴ�/�=�`O�Wi����u���)1Ξ�d�`O�½�3E�x\�����}�k�B�(��J����3н�W�]3�i����O�L������P��R���f�#`eSY�_�ߣC��@�0���Rҍ �0 DBe�� 7ڏJ��	�Nr��V�w}�����G=�����a�ҳyЀڒgIO]�ӝU;�Nr.�5#d��n+o�{r�8 �"|��	�����J�����$��)�+�fawh��sX|�7�n�w��{.��F/���c-�<
:�lYO���E�������=W�,D3 '�O�6�o?�&�s�/�t���d��־�'$�ٛu{���|;�P}�E�e�e�I:�������D��̙EL��m�̂*���s�N놵j�*^YL�Vaݭ|�L��?��Ki��I����t�C���-�N^\��-�ckU٠5�kS��M��5�p�a�A��ř����y�+x =��>��bI�e�O��]ױ5�
˺�@O�-3g/fv�����<�s4��4�����K��f0̖��i�g	.�T�ͬ����>�m�z��7��)0|$1�-@�S�ET�Uo��s�ˮ���|Ц���=�1ڷ�,Տ��Sx�ds�gk㴮����#5e^�N���߈q����{/:.��V����7{�ȡ��PUT�m��u��-"���z
ճ���q�xGgFy1ˇZ�x!�P�s�ARP�a�� ��#6׫��6s�����L�8�|�T�:cWF~5�g'$���2�	u�.�S���yn�o:�y{K3S1���%p�<��*�	�q��2k�;�c u����ې���+��u����l��}��?H�r�N�&JB���$�
��w5�8�|�Wc:0Sx���A,��=^��B ��
�����qX�>QiI�Ȥnj��Gn�P/��5�U�W��4��!Et3Ok�M��Tہ��	D���F~���kO�����`S�Z}�s����Rg��=I�w����A~��� D����4W�B�a��q�d�AX��
��2i[��*�r�-19bIdZ-X�*?[g�u~H��_f��R��FI�Y�����Y� `ˢ�q]��A+\�j0	�R2:&�{r����������8������Ҁ)�7[����nL�RI�Ԁa��_���9���c��T���D��g�z�#x�H�a�~t�M�_��6x*�*$�d�����~ �qU7����Ofi��\�Zwe����;��+,7�����&�t)�0�����9@o���a�F��o�q ��#�Z�%t*i�|vr}-4��hS��]�R�̀|Vj<C��#�áȏE�N�u��V��Q�̢f�B����^�<�=��e�W�D�?����f�[]�����v��l��#�)�S����Fr
0�e��� ����y�;i�Sl����i�WO��Tu��\)�=��!A���ĸ{�J�Q���Q��={Hw��p�׳؆��L+vB��� �k)Q��YKnl�>@�I�Q�/'XY_;YtA=��Q��m��TIZƕk��ߴA��b9��"h��ZXϣ������'���AB�
���0�x�����
�����ătW���Y&��Q .�9�[9qg�U��x2�%�a���)��J��i+�����h�ͣ��ȿ3u���)�5��x�-�	���օ֯u�~�M9Y9�[��{�x�o�������u�H���B�H��}�����M��ZQ��+hi�Eo8���a�sٍӱ�� ��;�gv�q�&�0�8�`�����!���l4��`�`��1�n��7kS\�X�e�Eg0(�ܨ[��Rw[��Mfm�gY�5ɸ{/˪�X	S��[��["+K!�j���<���N}�/&|T3�_w,�w���vS� ��Ư�(�:}��D�O"�VO'��OX�)����(�ab�g�
�%?k�lѮ+�g�����I��@ٗ�>"m��Ϛ]7��VS(>6�ަ��,Uu�`m�~��I�����o6&���Q�[j�)�z�)���|B��^��N�U�v�%�#S�9�9?iwe����}��)~hP ��8�<�����>*;������J�*c�6��%á�`�_0邒В��ӂ�Z�&���G)���n��h�5��G���+��!�z��.��ڬ[u (�^�Ca�F�s���倆)�s�.p�}�k5��spSB�lϞ��4���.p=[�2︑o���ޢz0�doo7�]髴u$���������L� ��P�hĴ�1!�h�6�Eӭ��B2��m������|ͅ�M?u���&�����qv��Ps����"������6A�#4��޺�Z�?�QvdZ�-��C˿dɥ��%�;��'yg�|�O��.�2Z������۠�U�?Yh�u4^=L_�e�H�����_-��<����k�KNU���)4�(.=�-,p7# �k��NX��8B�c-��p1�Ӎтb���1�P�:�%`g��,A �nV����8X0��>	�ٴ�Y��sO���y��'����A�C#ˆz<�Q t��|�ح/͢�N��0�M����f�5�MD�(�:�++R�e���4��z�	I��#�'�D�y���>�0uCi/�$�M���if$n���er��GVnH��31A�^����ۅ��nh�wfB8�_�g��=�ԧ�s��-0�qjY�?<�v@�2Ԇ�%��G�/�
a�/3�jjfsm�������9�6�?E�j���r/a�ۈ15�X��ܒ(/Ġ�(Z�k������#�?���;�c:�gnha7Bg��έ+,:L;&����F�۴����$g�/��!J��{O���p���MٹvE*}�`g�Nri���tEK8��Ia�
�	��td�o��oJ�6��v�����ڨח�~&jF�W�zbl���\>��̲|I|H�W�պ-�`�.�:�v�5�M[Ū_�H���G��RI*?�z�2w�j>�)> �-7<���]y�g��(_b�5�#��7�FG�8}�f�
,�wPE˩��!��a�ZF�8]x�9�7�R8�\���ݐ:@��z_A��c��]ɯ�^ˠb���������4J����{%�|��a�s�xS��>}k�H95o��8����~��~H�l�=�%ix�ѡ���w��bt����|\��������,�8݆�]��H��_q�T�&��Vp�(�	O���V/h�#��]Cjj����gH���\ћ�Y�t��&E�z�a�+t'�qA^�x$���-cT����&��k�]���:�8�!��	���#�8 ����'��&��rM*0�ي�i�E
&Լ�Cao6�K�hLw�P��M4k4~�8��1�B�k�i}Y!�`�ǘ ���沩tʱ�������z'��VY)y!w�c��\p�#��ے�b ��]��>1!z\��đ��t�1�+d�a<ŘSg���@�/6���`��l8٧b�����j+W�WlU�`�S���y�n�	Ƃ��Zx=��V�<�4ld�Ҧ��pEz�:�@��>�����<�Q���[��fK��{ݵ����dVn� ����5�Y�fW���Rt�~�Νe,
����2�9tY�WBoj���oW�qg8��d�"���*�gɣ'U��8��H1^��c ���"-ED�?����S�X�V����qߒi��Y�d�;�kƤK��/�[>)!t~Ҋ�Oɴ��n�p)%7��n2Q0N��CI�B'8t0VҪ���YK��]0wo�v���%&qf�|jq怈�f8ݕa)����9=�_�h]�M�B-z��/2!�s�<��I�{���~�fk�Y$��@^���Z޻�� f�_�
V�o���悹Qd�陦v�kH���u��(s����8sS(;dE�'`����'���b�ۂ��%�%�RM#Z�7��8�I����q��<�B�� ��ӈsъ�A�!����l���h����bUXc|�������Q���;""�@�k�0o	�9t�b2R��jBtS��
@�U��◬�Q��ϕ,ǹ��E�?��b~�I8��܎*cb�h��˟���PR$/���hY`�鳦�kQ��hR3����2��UI3!���_đByTh��P��3I9Z-!�m�o'=Ye'C�vV.��V���ɻ.&����;��Aa�����H�j8�/�V��>_�f�����;h-Sa�n�ʦ���(bX�\Z_���ô��B��J�l ��V���s]� ��%Lc���M�-�T;$;]N�3gY ��G�ȍxP���х��w�蘧J�]}���v���ң�{'��<���o�Ub&N�JB�3 �|7
M��u�M�����D�-�������蚈TO����Y	g_[��;�XQѧ%�;�t���~F��ݓ[��%VAu�v�-��ztpO=Ι�:��� azv���;�lpf�y�t}��q����̕����� ��?Q�GS0�{��}�\bB��O=��>�y%���F��
0n�
��-��ƃ��Sjz��b��D�����5�(f�w�8/6�ڊ��t��9�
!���Bszc�&�;[���v,��݉�	%ljX1(����ݻ�����W��6Q(d++��Y�1f�͹㵥N��AP�0YXi�%��uXp{�ѹ< �Խ�i�Q���#1�ԕ��2=�Ne|��-����6á��ak��7��L[1+�P��\o�:6����>�b�U�J�e^/m���Sq�%��11���eOo����FO�\�����]z��}��&}%7�g���
����.4�U�Ȳ����ݻa�|�����FD�*{̟md�m[���o0п�Nv��A�O4�^_�jTސ�?��; �wRl��ܻ��~���&XZb1��ϦS�����3\�k����|W$T4ū(��#iG1Ȉ��Bxط͇�8��6BwN��Y�?Ӫz�c�n�c_�����ΕF\�Bѣ�4,A�A/�f�{iEP�sA]�D�|oY��`B�N�.}��nQu<,��.EWY��K��T�:�e�e��[��]���/�B
�N�<R�A�{��b�����Q���U��ҏ�c���I�I��3�B������o�U�1"�ظ�57|̰�^�G����R5�5J�ɳ��0�O��#�v�T���f�`�Z��s]�W䛰�E���:����Q֋U����iW~ng�?y���c��.:ϕ��� �^��_�����;�D��?8")M��lnhI+iW��?�=oR�-�?�Eϲ>,����t��oR����-H���	}�d��)%V+�_�~��[61Kт}n��0f���BZ}V�����1=LЇ���=�[q%]����9� >k�5�͛�\��aR�{�6%��.3���[��X@�t��x�ٍϯA�y�#8�ų����e�i���x�Q'�&�����q���R�u�3���/z���G`�ڡ�Y�P(u����tG�퇆b���1��Ar	-���7`S��\|���4{6�ŕ��$��Ӫ��`���|@!�� �F����<���Z;�4�1\7�(6T��%�v�R�x\�1F��3��D��з�U%�^%�q���S!��j��L8�~H��5:�B����A�Ū)O��ʒEK�1�ә?������X�zJB����4�+�Kze�������o����\��ͫ�C�����/��M�%jaG;}O3���C�{X�M�[����v��:@���>�{�#]��Z��h���HM�p��|�A�ڬ�	j���X8������7��/f�rh�iViZ�����c��~wT!6waZ�d}�t�