��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� rā�SZ )����C.��&0C]�-��[�3�-���+��պݣ�k�J�vo`�A�����f����u�X���v�=�а���]Q�Wۿ�߸�=_Q�X����j>��Zw�K��SvX��ƥ.���#�����Z�0���#7{��\S$��@1I�QX~TQ�E��db����۰� ���>0�%�9�j汈��}��1� ��2���h�G��SeY�a���	'<x�p��k�H`�H�j^y�0�s�78+���ֳ�`�R3dW��_��{p[�?$�s0��#�zS�_��bH
�c�p�IL7]� |����Q�� ��Rr���=��E즕2%�����`�^��l�q-�]�p��jf��Ӽ-f%H���ȳ�>��+���M�71��4_�) 3�46h�rb�J�W� k�h~K0�>P$�_n)���5�r�j��W�J&޴o��$>��6��ŀ�;A~<6P��K�~��f��*I
�Z��}`q���ApC��n���g���3��-�іrO�mF���,�$��@�BI�q�}��Ȥ֐����î�䂧��@������U���vU������ �T#K@f�㯁����|95<@���+�-�)�����K���FI�k���*@�m&���
���ma1[�2�u�I�\�U�yu���o�|��2����;�W�W�}P�K>%5�'�8���׫=����k��,�t�M�0�8]q3���N�u��j�������ZJy�H�[`���W��b���-qJ��E����5q\bx�w>Ʀ��Ò���r�܂��%,��HഈdV�A^��k���ɖz�@�����K9w�5�i~���^��V���.���v핣����KXb��gt �K�1�<G��R�2�Yj�܃�)��T8յ�}𨁥�²� �rd�9�	8�y�mG��N��'xW�K�l�J��)zR-pć(�yN�7f����Q�GҪC@x�d|k�&�k�*�^M��F�jG�����{����R����_�v�wv��:c	\��������U&�}K���]��9�X�tReA�N�6��xVг�>'=D��ؕ^h���P���B"	�y%�-j	��^1y���t���]��x�BpVW�j��>vu��;�2 x)�ǹr3�k�k������2G��]��GҸ{�~L�ީ�X<M�?�$%^���ȂXY���&��u=sr,����ʢ��}r�c��Q�������,�;Ҫ#�MͥaޒP]��0_t;�.�q~�y�a��(׍��P�-G��b�y�_�q��f��'��ҷ./�������Bg�>�x��
�3g+16Ũ��!(��"�[Wt��_.�H����G�j����4Fy�+����B)/��7����1��"SK8��PQ��(#P�8\H x!sR܋�EÍ1��FT����-�F���E��hQ�������Ġ���i��E��A\ATq��|N��+�؝ה.9��e��Q�n������ ��C.���\�_���l��>#w�D��;��$p�" ������S���=�.6�8K�u�
��,��X$�mܴH�T&��-7���w��,�=,o��t�mN_Vi�H����a�w�	�g 7:���V1k��*�*�B��(�ּ�)m�|�,�]C��o��^�@Y�/���& �[�$�%f��)�.DQv�(a��t3$=���K:^�)i��X��� ��k�6K= �J�^J��f�MS�3J��V]T��׸�~��������V���ٲx�cf]:����H?���"�t)��o���Y��l6�L��{U���|ZI����@P8a����v��!�������)�Y5�D&|��+i6`�{��Q�y]�6"+> � ���TC��`p�]�9L�h��t6O���[j�!�K������WK�~�3�	Ag
7no|��eJ��j�+�p�B�p��`j�c[n69�{S���2�Vt�$�!�DNpH++�ՎJ]�i�{r��"�Y�
(]z)x�x�%4��=cq��.yҦ	�*����WwL�3����ss���R���č�S�:]Ƕ�Ua��^ʅN:tOC<��F�6*n)
L���^'��M�s���B.�6Z�Fx�,�f&bn� ����',��I����&�	}�̓�r��7o6UD��K�����j?�b�j3�s^\�Ye7?��O&���u��?T�7�vV&$PBP�3���|i�*?jŦ�!Q���"���!v6��K�2�'V���$H��� 9��?�Č�LXWHAД�ؐ�}p�b:��_Ys$\|�,7V��?˲�5�'~��V;��@Y<����6���k�w+���0��;�������I:�4~�����T���m��W�Ñ�$�e�dcW�+�\�M�|c��;@b9�ݒ�L|lo����Lj��Y5��� ��}'_��������u��ght,��"�M�Y�-�R��F.jw%���R%��<�ې��}*�0���T�����������Q}�������ģ�(���}�ְ6ĽufC�B䉥ĳ_>'�Xg�U5�"�C}�.m���IC���ir���]��Lk4�J�3�f!&�_T��N4RO��f��d5g�Z�K.{������u6L˿~J��P�5Ì���ǠtHw�$uNK[���rݫ��>��
Y��Eũx���݋��m?ND����JH�h׃�g[�>�
:�q2�e����u�#�7�JH�=jA����������⫅+��ijD�e�n|��I��<pn�^ ����_a_Ԕ����us�F&5��<MK4��&�*���h�J�pFf�Y�?G+l�9����]�h��Z��>[Ru�T�n�bC��_}�6mx�A)�\x8���Z/�;)j��<�>�#�6a�q�usEF�bͳ~��"_s��؂�����xsK�v�H�q&��%��F�0�70����(Ϝ�C?�2���M鯉B��Tt���#~ ^��~��Q��E+P��ڔ�f(��_H~�4�Wh�W�G��OW|8��o|h�yՇ9 �-}C���$ty˴,�I��朧�k�[^�����:��N&�o�嗪/e"�a��yX�`z�t�>�r��H+n`��0v�A�����0@���I�;���5�ēHIE @	:K���*�z�-qƋ��^���t�BK���wҊy)��I������
�5��C��F&hM�b	gr�
�^�����sb�x��j�G)��A{�#��7����2"���e��(��V!�aԐ4�C�����z%�9}Bћ�c��yX���$%�x�	[;��;*-�K[i��6��g�"����w6}r�L�qG��4Պ�	�W�N�D6i���2�!~��/�&�P��t	��3��x��86��>�%�q<��{�,��%�,�+Գ)"�
U��3�ǂK�h���e��{�CЄ�kjH�Z�}��/b�x����ƧL����Nr��F��t�P�����p 4Ũ ��%\�G�Z�H��pY��v�����0��A���������cVvћ����T,�j�Riρ]��+�T�t�.���R�#��m����9{����r����O*�aXP}��'�s2��B@�(������n��T��p��hw\��IX=�w�A�PjK���@�7>��Xa=R+,�cQ#*@���N�@�����P䳻��g4�ɾ�S�t��c2�MR�&;z���k�a��{���	�6�����I7�Zr ����\����,�SЗ�-";��G61�6K?k����E���Y���=�"�`��e�/�D�U�f�1#�kX���7fk��	�<�%)�ja�$4�*2�Q-��lI�}۠G���.UyڥXI=�@T�4��ax����Hl�yE��D�J��k�`�*xfu����f�*lO@������
Q�r�� 7:.�������K��ψ3�o$�L�h������	�����Y��mv9�s'�8=@z��2[# ��j��_J|