��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� rā�SZ )����C.��&0C]�-��[�3�-���+��պݣ�k�J�vo`�A�����f����u�X���v�=�а���]Q�Wۿ�߸�=_Q�X����j>��Zw�K��SvX��ƥ.���#�����Z�0���#7{��\S$��@1I�QX~TQ�E��db����۰� ���>0�%�9�j汈��}��1� ��2���h�G��SeY�a���	'<x�p��k�H`�H�j^y�0�s�78+���ֳ�`�R3dW��_��{p[�?$�s0��#�zS�_��bH
�c�p�IL7]� |����Q�� ��Rr���=��E즕2%�����`�^��l�q-�]�p��jf��Ӽ-f%H���ȳ�>��+���M�71��4_�) 3�46h�rb�J�W� k�h~K0�>P$�_n)���5�r�j��W�J&޴o��$>��6��ŀ�;A~<6P��K�~��f��*I
�Z��}`q���ApC��n���g���3��-�іrO�mF���,�$��@�BI�q�}��Ȥ֐����î�䂧��@������U���vU������ �T#K@f�㯁����|95<@���+�-�)�����K���FI�k���*@�m&���
���ma1[�2�u�I�\�U�yu���o�|��2����;�W�W�}P�K>%5�'�8���׫=����k��,�t�M�0�8]q3���N���GvZ�#z�HM���f5�����;�q��Pj����H�L�}��T7���z@�o	%�PFmy�lc�
)�8yIf�o���Z�"4��r���o�6˦��)��"�~���6��}�pY���]��
��K,�	���1D�̹�@��$���(_kk<| &���x,�u��Sm��Fģ	U��U9�k-��c�KU ��1$k�):h�����!�Έ>�l�B2A�V쉀�#� o�Aڐu�Q�%`��ܸ��cb.�����E��&�Ѯbz-V*�E���bnjۜb>W���z�<\UlA"���i��J��Xj݊���	p��k��1O:�$w%�C�\��H��U���Z�W��k�B�E��d��/���|�0�=o�g����/Z^����X@�N �Y*E�M��j��Ʒ�G��V��$��Qhw-J���,�B�����>�n�N9+���̍�)ТP��yw�~2�]�4�E�,��$&�_�������%�#P� M����PA��[�Z]�ϒ=!�ܠ��T�X�`2s��gq�D���&��%�?�Gy���4E��[4�͹��*�r�S�Q�����!P<�g����j�m2W|���i�:�?���_7��[�@k��v��I�������,��u�T�䷏Cë(��5<-�����8J���R�[{{l�Ijt�d�	0�:�K���}�� ��@W���D���&�b�kݿQ<
�d�dl�\aJ�n��En�V���pT���u!=��$�Z�
���Ѭ�!���w�*	k�����h}O��� ���� ���Q�����W0	�!�=Ť�A-˭P@S�� �f�3sc�D{o�nL�Fw\�&�ʮ��/�3{��U:S�%JowTc^��
/K��K"��6��;��)�jkxS0�+U!N)���0d|�b`�Q�?���HT��YMN,t�j�s ��c�M��<��e�l2��@C�dt�E^��)��NSz��I�<�h�|{vp�`�RL��w��h�VN���g��	�,�\�����<yu*��7�2`��q%��H��"b�U�
��V���Q�`ѥNN��,�''OR�ɯ�ql�b3��.`?�:�@����Yu�B��T�t�T�ʛ¯H޺�*t2�9�݋�B�����`�����șcd^��A�(M3��qji�j!;�K�zh>����:>GG���]�������a���m��<H����FzI����ݐL�����ф���N��������
 ���U�>2R���\���5:$�Nv2���c�f�JtxN-��e�Y�K����h9\d�T�S��e���/<��p���Z�s�����'c���k\0�,�Ma�F��DL)z7�`	n��{G�9����p��aǋ���1�a��1���J@y��q?�0J�� d����/�c �A��g����VY���e1�(#28��	{�R��Lf�b�ϔ�����+r~�n]�_H��8tk���[Ȝ��4�}@{�zV��|j�ژ�y���8y�R�>\_� ��S�3BH�_����W����d���q?O�	[�Y��Se�|��<��r�a�S��nG�
�ku<Pg�e���K���SD�,)=��8��θ�I��i�..��M�{I�������ua����ܒo<�T80ܯ���$��o���L�q���a�r�kZ2�,�K/�q�<�2㭠���̰���G�DIz���z�q�b�W�t@�x�,`�Riۧ����] ��ɐ�}Ie ��Nl ��dɱ�����,ԅ�{�ht񨑩Ԏ��,>+�j��@���ΰJ�? À�����D���$;Z�7�CP����\��2VX��^�y��Ɨ�-��V.
R%	s�_̨T3�7�3��]��ܒ�#Ũ����⯲a��I"�b��N��R���d���~(�Mh���I�N\��c��F$���[�k_A���$�븷���+
1�(��Jnv������˻ZL����~�����K�ؐ�s��<S�-���ͬ��^�[�ȑ�z{ �C�[�D�� ����tYu�t]��`#�WP����9"�[n1����:�;Gh������Y@i��&���S�pU�z?�8�bh�~����	���AA3;2"X�D,�l������-!c���4}rŧ��}�s� ?���^��F�������`��S�xp�p��5!Ho���|����&�����8�&�?�M�ug�]�6�����fP�����ϩ�^-��M��=L'�4�)�"�Ƃ	r�sI�@%w����ɝ���i�iE��-�d��m��\ivε�TK#H0�����.�s��� ֤�Nv�jƮ���/����L�p�}���G�s8z��񋚇��u�(,{�x4:�>?�!J�E�U�Q�P4�g㕲��+�Fgo�P��f�ondB��F�޻������غ�6�Q�~�����jy���i�Vo�4��@�{��s�VX,A��9~��X����
�30��2���ԧ�#�2^DӮu�HñZxUU�e=O&��Ol�ʑ
�1֜@�kN�#��N�Ml����P�^ ��A^�.�F��?���#z���7U�xԐ��|�<L�w����v����w@��H4F���}	kKA)�vm��I
�}#��ј�.3F*�0"�ZT�m��i��<vo9Q�,���>o|�"b�K�o����:Y:R�3��֑k2T[��ӝ���ފ���<��ػ� �$��М�<E#Fg��9�`�I@R<Iv^�m�Oּ�|���F���q	a�,[\����U;Wt�Fȏ�"f��q�'8H72�Ys�(b��
)��Œ��,�*���v �k�|��ǰF.ܘy8��N���b�v$�6����%��q=����Y`2�8'c8g�mqG��㙔��:L�r�4?�nuI���M����yZsGۻ��l,��H�����q(���n�5ۿG��H*']�������
[����5`�,5�O$����)A;yG0�'��A����p�������t�z}��(guJ�\�m�f_�b���I��ءL��}4��'�L�MX���;���X�lc�,��vZ��d�h��� )��T"����h�o�P�������1h,[�9�E�!p3�����?��,�j�m�|3a�n%��^3��zy�Z�i�)�0� !���}�މ�7��T��%�r]�\� �4�T�d��F��%hU�i/�u���WhN�K��ϧN���~?ż��aVqB&�=���P�]�;�ؘܵ;�F��FAI	W��r����P�N�Й"o$9��e���5���6�u�U��
���ۨ�є�;�t)V/bz��*���H�k�L�C�;�;��#`a�Ǆ��b���Q�-��9ǅ���|�%A�i�;��.����[ta���|�Ю���|��U7���5�^'����v���ù�\�:wu�ʆl*u^��h����g�h+%mK��a�к��0�ΐ��Ǆc�|Un����M �B��~𥘭V�&A����rz������b@u6-9k�9zx�� �Uz	��ol�����t�]M��[�'nx����\��Oe��!���j,X
+�U��{���ipb�"$?:Y)��Ȕ��7ĭ�6�\J擆�����T�����Y�N����2r�n�0�r=�J��̍���ޕ!�냄_!�hkQ��m]���G6U?�l��,�͉sb�a"�)��� )�)�%���}�t�2k� Z�oɳޒ����h�s��4��$�D����x�9z�%��r�k_g�ܢ܂�\P����[k�bb�ڹ��/+VG����y^�ty˫'��5�j�����ӳ\=$��� 6^;��0i>�5N���4l�E�� ę� �N�T�8k���	��|�R�r�ɎJ<7����b��Y q�����T��vz�7��wh�+���E�`z���g㓠�剌����7�
c�`25�F�Ej;������\d���H���!<|?')z�d�{`霫�3�
�A7�k�D�b+��s���
*��ԮT �H���T�۵�f���q�N,JE]�VX��%٭I�H}�o��8��]P��O�;_�:W,�yR9���$!1~kf4o�zC�^~��D/�V��]�RO�5w*DY���!�̤�+�!pg;��e4DBjh��1˼ϪTN��8�X�:��P+��Ң�7�r����� ��-�ьۅ�S��Ո_���&A��Z���W�g=n,y�t�Y̙Ο���ۥ��(��鲍z�]��C~�LHt5�V�C�:]���;R��n���8����ow�j�Ko5C����d1�%%�ydTT|��7*�u�r���oGd
|�J�MZ�i��V�7R����b�+��*a�O�h�w�<P�;�2ŉvg�%ah}�kl�ӝ;�-�K�}�Y�2k�ⷺS#�5R�hLsGj�ء�H����t�:�s'%u�7MO

DeK����V^N�{����Pr��fg���R�EU��@�B�+�K�U<n��-s{7�m�um�4�̗���+1ư0D�7�`����$���Ж�V��U��,p��ǁy�T�֠���Q��%1^'�����Ş$��@(c9��N�W恻���D�P^�%x?�c2�**�i�ٹ����@Ӱ_<$���b��a��:#��M���R�{q�{Q,J �;��M�z�bi-���Ų}��T6!���Jl����ah��~�������<�WVPlX��c�����F]`�.��n(v�Zq����σ��ސ��
/T�ǌ(h�\��~����Զ�ާY��V�|���O�\��$SI��M Fc 8RX��T.O����;h�u�KA��y�����zl0�#O��m�N֙������������$0?�9�tpn�K���T�,�����e�
�\'7������?^�}� �� L�����kj�����\���B2٪��p\`]�e�����rv����K)w��;2~��!��p�"�ӂ ]��T���y��!IY�>�A�]T� �i���"� x��� �Yq��I|��W�����D�i#b^�vaPU*]��V|��I��~��2����{F��(f��7I}KZ$�8�f�X�>\��ҫ�"d0�Å*�3��y�! W0S
O���o�,�
E�B�<4�^�x�-�g�����2��;=���Зׂh��4� ��s�T4U�3����
z����|��;�T�)rX�}�,aa�p�JG0$fJ���\� ����$��I��x$p���`��3�B��7�S���Fd��M��FF}�������Vs�¶�xp�FB��mk�
X�/ ����Z`�j���T+kG0�ﰓ��j�3�s�H}�,V��7%�P��9s:uڬ��\`l�݈�p���P�ܭE��z�$qǧ���ӗ ���{[,|��Kcg2�śfJ��XX��
��)1P�X�` }���5dᔤr��#�e�v��z��A�4O@;������x~]�����ڼ��"b�=)�;���VF�9�^U(������]H �"�7,��qp�,ޯ-�~9��ԕ�Շ5D���=L��G^;�"�>�V�/B�$����C+����,�ڿ����h�(�O}o�ɣ�*ӌ�a�����g}�[՝i�\�eȑ&I���:1��p-^u�L�l�'�9ehS5%~�r�T����|$(����{.�����^cH\U l��-���)��Ї;�~q?={z�E�
�1��R;mz�p��kxU=
A�@C�u
�t�5��,���Eۊ�]�c{EX�����BŘW4*U_2Q\�uS��4C�4�R@;���a�łl�-ͽGd�J�4Ռޥ�7�ә.";�0�&���Y�� ��R6o���<9���q�&]�e��˒T��4q=� Y�W������&sn���=�`+��Y�=�\����d���SLj��I�*E�1@�+uAv��(q'ڙMǁ_b�h�I6� !X�� �4�,���v��]{��	t��l�ם�����p��Lɢ�r0鉣�%�|>�C!]NOyA��LB�XМ�	s�0�@{e>_���zȵ5_�d`����:��M�����!��N�8S�e}�����y[���5u�a����jT���8&[�1�SϠ AULhPD�ù1*'��J	z�������_>����!-�R���Ip��z�����g��׺ؙ����0����Gn(m��O��ȹu�h$�QtGJ���9�k1�E�#.�/y�c'�
w�~+򒃃�jh�53�ޑz�/��nA}Έvd�D�P%'v�P�E� ׿����|s��d���&yw��2?w�Q"�;�]����3#�f�.	��T����gbǎX��ЛH�Bo�X����>�')B�G=Mp��E�cݹ� u���i��yd���H;	~2~2n��ve��Ե�)�CsE��}��ڱ����H�A*+Q(�A�î��ڼw�s�z�=���T	�lRH�_���\������:�����- ��9�TμN<�l�H���j���
OH��q�9����vh�2�����v���fѫ'���$3[�7r􃛦:�Z襳��C'���Mz���ю`I��v)E�&N�N�� �Q�@�/	�S�ɫE�Z�x���O3_$���,��3 �3$�<�~�(�ۙqipW(�o�+2Зw�@N�G�� �BAw���}2a�_��l����}d�'�?��8R�_$��8�W����w���.g�
61��|�"���_�M�C��Ig�6�$[ա�t��"ސ�/6~=�Ĝj[1X��H셯x��|�qB��]*U±��@UhK,�"K��;5X���E��Z��M\?r��ۼET�!l`�[���=fګ�L�u����"�;�y�������<������Y�E��1B9ʓ��	_ [%^����y��ܒ��[�U�c���T5�S6��@�+�گ� �թ�T�5�d�ԩ7�Û�}W�}Pj�!�"�h:]�v��w�0#K�\��w�6���!Ş�n����rR�R6h&���Ȼ�VJ%f�I��6��7��a����CT������~��8�j���Ůe��`����75�� ��"\
/��
�?v,�5�:��iL�c�[b�4r�Ʉ�e��Ι�kq͏�v.0�MԿ����V�x���-�eH҇�u7[���ˁ�N������&���Ψ�rWU'㻸�iI�b�����E�����%`VT�����},��U�p������S9��@���*����;*Y�5Y��غ��沦�R�V3p�袰ӯ����;j�'��V�Ѹ�`dt���s�]�s4�@Y6	$�z�8f?�Nf*��z���"N�� q3�
�w��M�l������>$��C%����Ӵ�Nk������~�竮د�f��s�������w�Y�WJ(
:�^
��X63�j�����\��R�CY�9�x�W��q�L��Q���GX�4�P��{-h�}����[�	{w�d��eF���߳Sx.8��k�c���\n���AKz����'�D��^�Y����W$���GN�R�-�w8�ͽ'Kh��@5��5y2<(���=6m$��@oN`��W��&�s���=2x*��\**U�>�HV�[u?�k��r��&0�7�=��;��%�8����Ǥ�8Jd������~��:��z"I0^�s�Z��c˲}RUR ��c��R�i���j����ݾ���S�F��ƈ������|IWV/�Slj�e5�Kee��W�v§z���|}&�{	��X��jH���<6(+�߃w@��.���wC�z�.��v�����&�z�͙��R%&?��ˋ�m& 16����7+��`'��Pz|/�� ���)]0`�U+E������w-&��;���o�&s���_-`_]�qw�
��6M=M���G�YK�7{��/��}V��G���'���)�~���X��w�a�N,�I�䒫B����Z��]����Ĝ"#�{<t���#��;���B��;FF���l�걲�z��@w/�	�{5Lf J��fqom��4q5��{��I�)}o Zè㤷0��B��%b���ud�r���5�.�JG�j�J�?}qƏ𓶖u�p����	@��+᠕��5fz���l������a竐5/�� ��'�=%�g��s�9�?�������oYKl.�lB��� ����z�.�l؏]oj���3V����Y�i��oP������Pߏ�9���w�C�p(I.ʁS��״��A��p�{r&���"Eخ�[�=w�c�y�I�
��痀3��s�V7uY�2�g�,��>��Or��+&k�fl:P)g���6��s��f��:���)��
�`��%�i��U�W�L;9��X1��bU��V��I��^ڃ�/Wh�Vl��H�Cz(H�N&��r-ݝO�͟ޡ'����V���	�<&F�}���4�O 8��V�Β@U$���U�"U�$�ek��o�Ѭdqw��`�w�"���:��H,W������/{�㰣�1[���h?�k7]��XU,���+�z����{�g��JӪ�!�3d"lg�΅�K�BS��~ˡ�����B�W���\�N��U�~ԵY���I1���/�t��j��d N̕�L�a�O�i�l\�����XG��j���b':jwdU�ҺC��	P�vQ��Dv�]ZY��^�8�@.�[�e�,����Oȫ�%�Z�6�vʍԿ��=H#�OV��n����q^�v�+�Fݑ>���;'>z�Þޯ^鷩�ۭ�"k7��%���7W���G��p��2"� ��� �'i�j"c�g��L�Y/5P0X�l@��a���Z�Q�6&<!��a��o0�׋����)YX�A{�g��ӑ�o����m^k���	S�_���B���/:ӏ�8�$UJA�(�
�tm�i��z�-w��΍-J6*��wM�{�}���6��&g�)��D
��Ꮮ��J>l�ȏV��