��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� rā�SZ )����C.��&0C]�-��[�3�-���+��պݣ�k�J�vo`�A�����f����u�X���v�=�а���]Q�Wۿ�߸�=_Q�X����j>��Zw�K��SvX��ƥ.���#�����Z�0���#7{��\S$��@1I�QX~TQ�E��db����۰� ���>0�%�9�j汈��}��1� ��2���h�G��SeY�a���	'<x�p��k�H`�H�j^y�0�s�78+���ֳ�`�R3dW��_��{p[�?$�s0��#�zS�_��bH
�c�p�IL7]� |����Q�� ��Rr���=��E즕2%�����`�^��l�q-�]�p��jf��Ӽ-f%H���ȳ�>��+���M�71��4_�) 3�46h�rb�J�W� k�h~K0�>P$�_n)���5�r�j��W�J&޴o��$>��6��ŀ�;A~<6P��K�~��f��*I
�Z��}`q���ApC��n���g���3��-�іrO�mF���,�$��@�BI�q�}��Ȥ֐����î�䂧��@������U���vU������ �T#K@f�㯁����|95<@���+�-�)�����K���FI�k���*@�m&���
���ma1[�2�u�I�\�U�yu���o�|��2����;�W�W�}P�K>%5�'�8���׫=����k��,�t�M�0�8]q3���N�u��j�������ZJy�H�[`���W��b���-qJ��E����5q\bx�2Tc�eyK�US��d�n���
јl�E{���3��4�X�jy�b�G���Q��P�`�����;Qm����E�g��j��hp5���1�]�"�4�����Z�v~��ާ���="��J͕9�CGӕ�Q�,Z�B����icek���6��f��V*��Hڿ�~U����6��`������Ќzw�&��B1i|t��pw�vx>�q���|XW`���жF暛�y�K1q<WQjE(;�/2�ğ��7t��>���~���l׍�� rq���U�x���f�������f�B>b����G��Q#�u�	k�����:�#�ʅ��}�u���k�$J���Z��ojIY���|��M���<���ip��H��^N��'�Mvp%s�yN�/�q��uSl;Y8����Ӫ��%�~1ÁK��Z+�|t�&�o۪#-�oE��n���)��e1�uIU�n$Z"����E��+yπ|6`���D�nu�>��s�T����,�
�u�x�u�; L�~�׌5�IeQ*����f���m-�)��3�h��H ���inQ@�C�2��vE���;yp)q�r�����跨Hs.��_����j������#�F�A�O��/_|+�+B
����������D�Qu�lI
	:���%^�2�xQÛo]Y���ũ�����`�X���X��6Va�n)�?�g\����Ʌ�z&'?�7$K�i5��PٌG�r}<Nr!��Xύ����l�ޒ��p��ג�h�l��k���p�޹`�5��M���|�C�������2wXح!}�B:gg&��x#�O(���F �j�҂���T���x�Du���h̻mIH�C҇PۯȑՙSAIY��`"���d�dU<K����踼~�Ѥ�LmyW����*5� o�vR��`Q�6%&w�<W��],���n�gi')�o�~�	q�b.�Z���f�)�M���'�'��zJr����Xc�e�Y�h�w/8�w�k<�B�ҁ��^�����$����<���EgTpI&�+ϲ7��7�[���{�0���jü���t°m�#��/�>©��ο~��zt�>��a�3�.�)��Ki'�V�2O��(��~���aE������<�[���>���"�i|k���,tO�'i���^l�I	L�M�	J���|l5I͐�{�Ez9��jᨧ::��ˇT9)9F���h�VQH����@Ԙ��B>~�c%+�I(c���pab0��E�K��l�:!�ޣ>+�9�B���v��u(�����@m"^�o���f8aw��J��<ޅg�!w�;���[��h��FOЧdx��Ov�=�Ё1�~��K�`����蓟ૣ��u+��U-��S_�v)����5���,-(�@7�ep�\o��l&ݭr��X�MIp�`�^)0�k�B�k�fK�p�]![���wȾ�J�;LJ9'�QhG@q����8�f�A���mΦy��1p 7�ZL�*2&	) �ܕ�_�����L`W�~}�6*����/��]\̀=�ĭ��^-?�㌑v��(�w�B:Fm�L���.�?�	�.�&Q�)2$�}���� ����X����rV�2��Q��������E�D��5��9��3��n kp'� Q������:������$q��_�=<A��߽\���h(%�N������4,s�V�pg�wb��z�<(��hB�7jFXGL��\6���9)�g
C�J�ue՟�`�1إ�e�ַ�G�u�$�L 8����l�ū��]�f�P�IG�iV��[M�g�˳^�����bU��FY6>�Ou����AO�m�]	�GD @��h�┋]��,Td�>�w�9#��"R:��;Y\)VͿ���H&/��!�"Mi$3���,��\�t���)�/�;ӇF�ltr�V����^�0�Np �N҅]���z���ahUg�~�Z)�<9>�!����G3)�D$|X4 _*'��q��r�$(H��3ǁI �R���C��f�9xC��6x����}�+��&�u���ܖ,�P�0�Ե]�'�J��u�$`E��+I��^�u�Om1���5�bK"�A�qKAf$��Ƕ~
;|Z������h�fΣ��TP�%�∀����|[�8o��Y�aO4�#<�k�G��GN�KEw��6�ԉ� �7
ud��7qR���ɘ@b��T2���v�!��2�#oQӉ���:gF�< ���[/)�ZO#}���!W�_�\<P�
����o��h��v����� E�=�
�U��cĵ	x�TA����x���]T�$_�fU�є�I�<:��w�.����))�E&S5 �a���q��j�)�g-J"�(�뙷愒��dEi�>����K͎���rP[~���9,;��R�;oIr�d�7Q[��n�Kee�Eh�Y�ݜ�|!�KZN�y'����Xn�
����/��,嬤�J�L��?���g��J�ֱӕ�7�j#{�W_���`Cs�
f������Q $R�NZ�'��+%m�xz��r����N��
%}��l��KNu��\��(vz%�ʈ��r������q�=W�{���w���|�I����^2�(${rWv��q�����_��W	�ᠬjH�9��g����q����$(�f�
� �K�y���c C��6q��i߫ӛr 5��Z����VË���Ԋo�����kщ��l����擪<t�^�b>ʣ��MӏIE�V)~Z�C	����1]�4M�v]��`b�Ҁ^mB��<�
`{����.����Z�S�;Ȱ�<J����3��y�[r���
�|�\T*vcRv���j��agWGE$Ҧ�p���q(������A�l�k\咄�
��t"�L�u�!GW/	զ�>dQk�� #>�����>>mw)!�M�S��HLZ@�:.�7�u%���ճ�C�_��{-LZܫ�/w%E��9����wr��o�p�膇��-��x�G	�w�����F�3N���Dv�U�u���9V��*�U.�A,����	�����D5R�
_��Z2�
��]uxo��Z7s��1[w8�|@���c��J;zz��!ȃ�h�k#+�E�%�R&��;���sƗ�fi��S�:��c�B�1�?;�Vw�|~���R�I@�k�ë<�;���*A<��������#�"� )Q.f�:eS�S�.#�D�X畗Q�:�]����
'q�]��i^�C�1s�����gz�3��~w6TZⰳ�1�00S���"f�p3T�8��A�)8��]'O�GQp;tc�*$JMm�V����n��h� �^�����g��;����2��룧2W)�JMG��H�7?l�y\�{L�Ibt��d�ʐmsp5����I1)�l�j�aO��b����{��k�"��lg�wz'����16j���
;;�	��SLX���c�21�̲�զ��V�P4�O���jo5|�jp0����#�]$��ZF�����T��C	��D�~��Z��n��1v��P���PO�YCG),�c�S �(Z[�\<F��	�D�P���Z��z,�oM�S�������=uo��a�r��A �J��*tFOc�W��Cce_�X��K��ܲ�HQ�6���3bm,^�xw�?��dg,"�"�
+������߉S#�8A�p�n���2;��l��-,�V�u�\e�I��D�g%s���k�=]�v����"�ɭ�e����D��]F}r�0o�j1��3����+��*��|�_��] $���L.���˃��.G&2ړ���8E���=H���QF�T>1��6�Gꛖ��-g!õ��7����&c���ɂ���g��^8��=㪳y�ӂą���@1)J"#<����7��}9Y�ı�O��>n�g��y�1�y�z�:�oݿ����ܩ�;.�D� ��i�xY��3`v�~����W԰v."��j2����8�1YDX7�T�!Q��WN��G��V�&.���Be�?�2�)����|�a���=���]��t\��,2�a`�\������3�5"(���}��+ݶ�R8�	�ޝ�X��d��t�.'��J?	�0TS���U2~<��zA��NuMVu����B�=�I�tP��i�+�06V�n'�����El�O�P٪
|�qP���W����Jsr�c��9ƛ+�׼Zq!��8D��c��y���+�����ֲڦ�]�*=������W�v¦�a%ǌ$�v�:���q���6c����#D��oZJM����^����Ȥ{Q*e��ɭ>i��g�����˹h�Q�f���lbO!.�寋���-_6S�wgS��"�8�H�5+�v1�Q�S��h�>�߄�����%������zgM��X'�b�ĵbNr�$��rE�{����c�Ɗ~��tͺ�V��l8�*)7��z(��N2��0p9�g߄7Q?;�yJ����b���88�T$�G�"�ʟ� �t��&��.R�]TN�
V�ش����G�I�#�\�+��U�4��_Y���*P��\]�C��Ls�-*~�oL����ɷ�gۜ �	�E�pX�B_ �{��;b_/Uj|��U�\�C���rd� `�Wx�VF�\��u�Lڠ��s1���Kv�A%�6N��ϛ���]�f�=j�
0�"���_&R4I«����3���*8	 n'�<�V�ow�� Fo;�/�]������%k��x�����������hH4��s�GZO���g�p�u( ������9<fS#�;v�I���_r>��g����ʇ?��|>FA�t5U���ݯj�����A��cb`�w����_A)��\8�'�ֳ�Jn��0�7��]�A"&10�/�����z��e=4�?ϯ�1�L�
��Ll��c���϶��îv�-j,�?�E���I���X,m��'��15��j�]��a���G��y��E,7����qd4���Q4�����&�<���a�\j�#>�9��cBM�@AW��샌:-PL�BwU��GP���̀����i*L���ʬ� �,"�$�9���%oo�K�4Z0�7�!���$b55Ȓ�wBK ����_0!�N�8��՟9��E�/tM�qWc(WB�4 �-zOvb��%��tdq	��״1zp?z�u��*��+%���ط3��O�����Q���p5C� }
:~k�eQP��K�>�>˱�ny7�����%������fGOW�Xo]���@�r]�mo���"E%r��Hi�5���1�s�?�xa%D�d/-�wIc�F#�Ø3�fr^���0�	w�ɀ.� }/���4'$�G��9���I5bO��j�������$½���"�*�&�K?�)3�8|������I�����fRF� �Bsҽ�Vsն�3��叵D7�=����,>U�}�0.�9~� -���+G����i�	��,�L�^Y�̔�h
/5痧�>,��w�'�#���v���ꉬ?�h���XL�Ӛ��!�|U�F�\٤P`N��|�]jPd���b&�{QzgǗ�͙�9��\�(I/��W[<O_rx,3|��&�k9x�	�JI.|Ws�;O�d���C���֥��j�#�;<|a���&[�pP�5�"?m~���)��+�TJ�DszE&�^�}�7��Ez"�v�S���6\��giسJ���Q�����x�w'}YZa�Ϭ�|��$���򣡵mdC`��(h��T�ũ���ս�|�t� =������$`��oT:0��k�s�j`Fw���;(�6��70f[�9)_#b>����=�|�y�fd�,	e�_
&Z*N���@X#P�/�U{l����j+��dРR@�PhB뼛 /��eT:�g���#� W�2Ni���#L�]�7�eM�l��ԾJO���������{M�Q�ƾ\��i�y&���bu��s�W�H�J��܈%E5�����r�Y&�ɪ@��I}
l`3�\}��j�N�HT�����
{�8�L�W�e��PY\n�K8���s�=���	�pC+
��%f�.V�x>�n:�5��Z���F���bwD�¥�~0�-2A�p5	�f-C?��U���a@�޾�Ɋi�w<CȬ��������P;���YQ��
��
A��0�-&���a�ծ5�IH�o�k�!]��@��~��XG�\��e�k�v�0��q��p���q�Y_i�k�?��}-��g���a�~��#{#R���P�w0{�� 8	�=�50)�c�����`�'��Q7é��:�ə."{�? �sK;��@/����l�ⓓM8̣Q��#��u:�~�mI��&��'Į�e��	b�:KF�\R9`�����0���j�<�{���CO�BP�o�"@e���#Oݨ���	��_E9�?y
ř����c���'�2z>�Z)1k4��i���󵈵F����$���G.�$��m����sC��PB[w�+F�Ϣ�צ�����Q˗ �*%O��Fɟ��Uc(��"k�=0� ������%լr�N�5����%�Hs`7�u=�%@G�*L_ $�,6�~�����
�9�:���`%�1^'��x�A9� �%����@����~5�y$Ġ�����&�h�o6 �A�ۻ�� ��]�>{}��9���������ʪ>�ZYs H~��Sv�Y���� �b,��A��Kk[�|4�{\n���Ҡj<��o��}�� ���]��qe�_���4�
�u�`��6��0�E��4Ǥ�J�/g�z�	\r1\���E|��Y/A�'���f�W����F!�8&�q����p�p��h�'�}���u�y�����ģ�^(`Vf�~gy�Ar�D9��a����GL9
��,���t�9O3��P��=ZR`q*�H�s�&��DW�|5���D*��c�~�S9��LO����� ES�c���J�<c�t�]Z�a��6I;�/����]��$㯀��zƆO�W-��~�!^��S�Hs����S!Qd���I�,��o6x�pV-��EK�#�`�w��� ��5�ֽz�\H>+ ػ@���b�J|l)���K�����L����~��苩���a��2:-w���U������F�ճ�$���2�yDp�v�IZ�	J�Rƿ��"�HN�9��x3_wb�4��o��yT�.��I���I����AdAE���=F�R��ɝ��,�˱��@���`X���@���N�O�4G؀[��#"�8�k�}ܘ�Z��ȷ�.��v1@tv�c�������+�+�I"l��A��n"&]��M��d��j��h����VW`��'��GL�.
����(����� �?���z�����;�wB��,�i�j4W������o3����k�¡�����8�����dT4��ʔg�6��+z�}��D��E(�Ow�rY�t�@hb��$:�_V"C Z&���s�� ��|��'�۲���y| �@�]AJi�5$�G���d���Pϡ����6R�I`|�/+:�a�Oi��q/A�����aF�[���׈o�,[���xr��Jv�/�<����Ol��5vA6|�l9h����ٙ�a�d��5 7i=8DI�s�pv�%�I~�R��1)�i��lį4��`P��ux�ņ�����.�<�x� wHI�˥�gѓ���J2+<q�(*P������C��S�4nv�Jr�}Ya��H�c���ȥ��R��C�k{A� d䢶�`�l���ߣ^���{����`��N#�m�>�����X��8�sp�������GO��g�nk�9��|g���M�k/�xos�����u�l�;�K��oޅL�l������9���ަ�/��D
��s#�eaZ���8gr��A�0�Q�+��Y=d�C�/�V/�)�V�f|>aaH,r��`*�
`��W��G�q�؊�wk>mqI�CJ���)SW	
%��g����o6e�X��ZU��H��K�+�7��{,��1�i;���UF�)MP�	���􂳸풙}f!mx��Jv��G�L���]�5s�x�U�X��ݦ�3񍾐$Жw�s���`n�a�Ҷ��x��(����݌���Q�p=�{��r�Cmd���(,-�Dֹ3�i�+�wSc�/��L4dt�
�5�}��h�d-=����h�8�Z�r�Ѷ
i��w�\*�{'�3���P�����	�\�~�}+p�����G&"��+N��an�u~Z���$"�pVռ	]P�=��U��v7��h���)�}hO�I㰅����5®4(Au��b�n_1�����I����ɀ��I��}��	���t�呵��Jަ�@xwP��z"��
�����l/ō���^�)�4�V^7�ɪfn��a;R����K&�6}��;oƎ����P�燾<���J�=[����([�\a�{�bw�30����۽��r*m����0 �g�T�U@'�tU�8�x�>�ub��;�1�W�]��!�-����Z͸⽎�uB�	��ʦ���kC`Ӓgy��9�O��{s�_��M��J��WK��x �;��u����{�J_�]�*�BW(zpc��K%����k\����/����N嗤M�cň�ppS����x�Z����TwV���7~ژrg��b�\U=E�+�͏�ǈ���	)�1�1��D/=�Y4C��{P�\K��=�<�����ߐ����h�*�1)�P�j(���:����������Ă�vC�?~b����1��Z��B-�{����Ǵ4D�i��'�iqL%A��Eg7�z!�S=LMR�~S��׳� �>�ڦt¢��7Z@y{����Tzڠw�����[� P��8:Ƚ1-�*�r̾�t�E6�tA�ԣ-�/tYP
qu�	F��D=s{�,D<1儵��*�M&_�E��"���tL�����T-�{q�5`��k�����f����F���D�Gwi�4��x϶6���x��Y�u��z����&6y\�j�[�ч����6ڌ\�t�|^��.�B�q�6�B>��қ�7��&�k2���J��a�2u�i���6e��m���0�mF�̡٢+�qB��M�!P7LT�+������3"�LR4w_F�\A0�"��ᤷ��p�H�F6���
�P����#rV�7u��ݦث�ͧ�$�|qNF
1��xl�-�x��mI=��br��i�:�ܢw��>��<�I5��k��F����k��-�?����oc��L�7��c�a�:��Y\V�هF �.k����"�p�D��jd7g Co��<��2���~�{�c���҄�%�?_uL�ӥ>)p�72�J`qՒ���S�5���P�7u�x����,q�Qu�h�60�ÆE��!uI[љ��<Tȷ��Mӡ���zd{�仸��p��Eq����D��\���r}��P�*T�K#�x��Ha�9�X�b�����3s��3��g�)�4{P����1u�]���"�[Q[f�Bp�S�ь�u�%..�QrC�6y����@�\R��V�1�/(�����k@ܮ��1Nʨ�Fx��D>����`iH����E��m�'hd�m��_��p�I=+L�<��ei��|�0-)8v��]��!D���R�hUx�}鶇ݬ�M�b�}c�������j�ي�yU�G���&����H�No(���:f�k���=<m^í���S��}3��-�v�0�ډzI+H��	JJ3���A7YD
F���ǙÏU�yѶ���7ou�8M������H�h����mZ��2^�X��on��;�kQB�]���p4&�O̟#�����|Mҭ�9���3(w��E6�}7Nx��Ls�K�>.R���6x���"�A���eE�����C�Vh15s��-��dv��O�M�U�V�b5 \�%�_0El��k3��Cܺ9,�4=@�i���]bNFW��B���K�%��;�6t5��o<�<2d���9�`~/q��kc2
V1'��M���/ݞ�����6f�A���<R�R����4��D�ެsN�xG��:�,�����7�|��" $h��q>	�W��gr�)���g����&�߿���;S����}�<�0�x�]}"�ʥK�G�1"]�����LF	@I��R��^}j�ṜoM	��h��`��Of��j�k�UZ�`���"U�<"����ᬔ���D�����֙�͈�;�\���+!6N��F!�(�]�����L�#��*����/��Ou��޻��0Q]̟S
�Ԓ��$V�>:Q�}ӆ�Vu5Ɠ��ٔ�j~�&��
I���Q�@g"Y
����Z��_�=Q�-4���|�Un߈Ϳ�5�4⦷�׎�����p껓�W	{B�1��K+������L�E����XO�����XN7�M���b/�S3/T~�v�XQ�X�5�'���C����L�=�z��R�ݠ���]%�ϴ'3P�!nΆ���Fc���t�hݴ�}0�k9�6@FB�{���ә9�% �]22����%I��H�5nv�-�cu�uH���x~��j"����Q�B�C$`��¹�$�A����D#�w�g�	g7�G,�����/���SJv�Dz�BU$�b��Kx	A�x2�;�kt֨��Ga�Z��u��ـ�+ؓ)��*Z/=�"3\ƍ�!�RU5���LiG����F[����>l�:fQ���!bg[�5�C��~�J,�`,�OS���@�H�=2[�yR+��B2K�^Hy�΢�:>��:�I�����v���A�e�,:˄�����=�x̄�0��!�57sӄl���10A�8@�!�O�b�,̞���/��]��37RaVR����ɀ�3��vL�����C�5��8הTN����& �r���7�PPT�H�bih����u��ve[G�I�A�H�)#E0�:�bFb%T9��[��������\n�2o�P��Xb�)�'.�e�j
�
�o
��:|�)�ǕZ
�P�ݟ�q�à|/���Q\�:�b�Su��{B�H� ��M%�Pe%��z��EXD�����Jkw�'G�lw�)��`-�Io��e�F`�m ��v��=�ൖ:�̸��DB-~)$K�}��p�@	���+Y�<��r�,�g>���n~EHq����ʖ��aZ���/�%���)i���������R���]&�r4���/�qk͌;X"�����f0� ðv}'9�!��}�:�-�0��i1�Q����-?Г�̲��I|;�Ge�Qh`�?��O�w>к{3��˔�K��ɐ�Y>��d��AT�U��������J���3�����q�¢�?�:���J��2�޶"�����A���J� �"H?��3�3{+ÀM��0�ǔ�G,�Ι�%*Ә;5���ҭC��[�=��� ���+�n�g�BA	��� �Z_��z����ҁl��,���~��:;$�XŹW\�To뻺@�i@]�k4r�RYks�0�y�ʊ�9�w�:�9�����Ø�rZ���8sn;�_A��1���܁�������BG7�q�W�93wz�}��dP�E�eUל�����<F`Y��U�'�No���s,oa��p���d'�y�����5�nA�)^���9�y` ���7�k�+�%�iS���{�QɭW���V&,;���3Ơ#k�	*
��6�,l�V"�>I^kx��+I��7�ga�	'(�jS8z�f:Hcc������'4ܿ�w�k�;W#W�h���2s8˙.�u.���|d6g?���O�-�PbO���8��P=]�V�~JX
@��������8'8�J�O 
��q��1nJ�w�d�����i���j���X�s�j����#-��������r5*����U�m]y��t$�&�c�3�D"Go��<EǬ�A-:���_g0���=c�H�g�DP�e��5��F��UJPz�M����/D�|EHǐ�W;:i��ڰ�����Xt[�Ym%]��׫J�+��%ird?96�{��lt�B��6/W:²`1� ����~�w�1|�+�)Kq����zz�`���"��u�J�(x�7J	3�6���hD[ٌ��{�:G��1^�����	�I��e���g$B�T64&!ђ����� 鶞ݛ�(�{�=���`q���e��>LE�Gύs��L�P$,vV6�����ͱͨ	`�K-�҃��N��liD��n&6;K��±*�V��F�`�Q�xjocq�^�g�2u�/�z�����ȿu=��`yfR[e�#�ڀ�`m�b�c���U2C�ÕW�G!��Z�6x�S>(�/N샌�����h�$-s"��U�YEZ���p3:����<�Kʃ?�Ұ�&�܎ٮ���:7�WL�H9Z.x:+�G��ۉ,�Rpj�r:4�.��|�8DKE̚������(�RM�/��mHlDN�.�:�ϙ-����0UF�����������y��;Դ�Er��0���!��x�*�K"�d�fϜF��h�S4~�Ul���Z�`��3��*�X �&�c:U�ė���('[�G��{dAW$�=��)a۵��LC�s��?
Ԅ�9��/�/�84��9����H��f&>�L=�Jt��+�mDf�9�b��^Ѕ�L�M�+F�to�g<z1�C/I��Fەc�1���~
�;m�Uu���9a6˽l��,�����z63B9%�Q�{	�h��b�~�� %�_7�)�_�7*[�I�R�Xx9-����C�,�⩗R�1�HDe��x,м�\�4s���+�9I4<HE���Gj���=W:ܬ�Z�$����s��2�R�K����Z�f��p�M��f-�6��:�X���L�+~M�hn�8[k��I� *�ͻ�������L4)��a�P2}���n�\Hq�6�LqƓ��R�q�������YL�{�̎�#����̢�a�m�k�cm���-�5��K��r,��WV\L�������z�!HR��"�
qnb,a��s��ۜ���U@�p��A�� 
^�l�idY�u64<�6Vl�/m��Ztl���R�9]�D��t嬼���/1Du�20O����a���{�
(�=�"�Q+s�B��A��=tB_o�_�A ���N�>U����h~���p+��8[T��횏� ���j�b�EM��I����:������%�N�(܋bUҊ��=r�ɛ�V����<�V�<��0�ZN��+�w
X�2bl���%��Nb��Ҵ��l��>rp�N��Vy����1���K�^�s|�*h�r0޽�R� ������B��u����*�e���H#|�̎Wp\p+�ǲ4�ʾ� ;T��*�{�S��9��x�0]�t��� ?ND����˽�VA
�P[�$z�o��cR��{s���㫧7��5a��cT@������M
�Us7���ʉ������]͟��/=n�1�)>�`�?�{i��Q��TS�i�\gJ�-��\!�$ڦ�>l�|�5�j�-Q����c�����C�}��8��h�?�?pr����v��� �:Cy�7�
B���kU>=��,�p�0 ٴ>fJ�SI?)rB�j6�Oo
6������͚������8���z6���.&�����t���T�o�[c�|����Tu��]�h2�{��w&,���t���*t�d
Ԣk���_�%~O'�7^ghR��Kp��7�t��K�l��5��S�}�H�k�� u^,����8��M�V}'��d�N���&��������	o���˝����E�d���XW:[�O(Y\���3*�I�V�c�rE%)v��),𶴚��s@��u��J�h�4y�$ZѡR�a�����4� ��{"oV�C]l��Q�8�lZ�y�k���c����wW��³!�P�+ia�j����<���6�@N�ϰqm��`S3��̫�M���	2�Hf����K$�ܸ���o�r��n��a}����HD��=�=�dl�_��0~_������{C�3i�~T��"��R^c��Ba^B�����zƈ�WbEbmf�����Ф��X�g2n��y�$ɨE!L��1����8�m�K���o�ӡ]+/��-��I;�^�W���+�ᒈ�[�����z���Qw�3%|V$?�㉃1��x��Z�^��-$�=��$4����U�;�M#���mʴ�`ω�*�����E�a{����C��Å�܆3 6OAN-�{s��Ih2q���D�
�/���.Rc(<���=�R�v�-�cS�m
���z��MU��J�,���AR�*�鼴����3������u�~��l�-�O��߿x�je��ĥf��+�g�%�v�:俪�
��#�)�'EZˬ��V�O<�,�L�JV)�8P�Q� �k��%@k3Ÿ��-ӂ�X�BB_�)8����H����mXHR���h�Pn���.���@�p�2��/3Ph�+������$(�k$`��F�L��_�ƫ4xO��>�%�N�nI�!����<�>7�3,�iOI�(�7�ݐ�n����VΊ�z���'6��U� ��� Ӈ�QܡMI�,D� q�e��DU�
�>vI�c+�0�2
��	�0`�T�n6����m��k��+a���3A�`�t�*�(l�o�R��E��iT� U0­�EXU袸+�+(�G��3�[a�c7�[4�!?W�,Ce��sY�g?">�P$�T�1F{�|��f�;�HN/d��w��D�p���"d��8�8<U�k�ZO�P�n�-����N�i'��	�є�6�m�6���w����ٗ$
��$B"�l�'#~��b�z�����e��E�_3��� >;j��:=�Ƹ�?���0T��������]�d�S�#	+_g �C��L�٩��i3%٫��d���r�"FI�w,����U��V&�g�.�e"�q��5���'�ԕ�zͲ��f� )c�i�F���2�Dԉ�iz�U�+�$��ymo��N�T�N9���j]�?/Ե�|r�GC�]� >&�~@�c�b5��P+�㚰�-��P*x���[��b��@<�a�{���:�C��,���k����x4�Q����F�b��E�fW3�]�]Ζ�}ϑ4g�BMgWnQ�Ϣ<��mq�YWO�5���U��`_�ɓ1"�pp��y'��;l��)�w�����r�:�eU�,�K�h�Ǣl�Q��J���oD���E9]��m,����|f���-�B����i��.��TSTT�f
/����������[F{A,@8�ri�o���I����WOא���Z�2
��9�I�����Gp�����ڋe�b�[�}�$����aLN���+��썲?7§@�M���D'z���R�`O�	��"����'��\��[�2��g��L��z6������hǩG���lRګ�`e{�lĊ����@��jP�P�D�=�JD��erʋ��v>[���[KR��8'���.Y`��{�M�l:n����I���q e��ۥؾ��B�{���<��Z��Ə{�I��a&(N̬՞���E(Y��L�b��Q�r�B#����7	:M�l�o�j~�L.za�o&�����9���1(�xQxω�T(D��O���҆�����5�g/�d�0Ձ[G��l�6�]�Zpa��[(̞y���u�B����Y�݄��։pEu���H�1��k̑��o�l��@���|@=�y��{-7���4.xn�5�4���X9+��lat��}E�_Q4�d%�d˩��A�c=y��$:�T��q/_�D�q��h{�}��S͜�xy>ٳ���#;�R��DU빿���:�an�k) �*�˂�Z������A�"�W��%���}Voee·�͖�(�0-���
�̬8��"(�-%��ii��=�s����U&�\"1Ռ�T [9��}�!��|�W��<,ۢ���Mf���v�k^��>S+�
��3����EE�� �Vs[��+
,�yr��j��z#�k�E��1q���e7����I�j��'B#��d�eԷ��ݢ=�,`�yy=�a�� �E#9�ʇ��ց�����e�[cX��oL�0�0��PV!����g��l)J���A���g�KއыP)����D���<?�uԑ8��ؠ� @ۘ ���9� ����RL����J�S������ĢQ���{ա�LHT+wQ�Ѷ�w�P��y���@����w[����0є�p�!4��d�-�o�I<�D_�W}d�t%��*�(�a�ioMn�*AƷ�b��Sy3�๯��g����<��@S<�V3�5�h���N�Cg.�בa�s��%�-������Z��s�Ӧ<�h#�Ưnl�_FL�Hjz�6�F�H$�l>Ƅ��'7���}6������	�@���3�A���uo�%( �[�o��p����Oa��mo����pA�rm�o((��8�'><Ώ��^b��ؓ�n�D_J�J=W�@�Ȓ�a����[�Obd�!+}��&]u������-��˯d�U���Ԋ�xPȶ0��+l̔ޥ�a��5CQ��0^6�^E{�L(FO�U�\�|�*�����f�)g;x�J/{���	1φQ�i�7��hf$sԅF�m�q? ������L��6���D��2V77Wu���HJ=	$VU �l���s���i�Ԍ?��_��e�0L�M  ���Ck�:&�\kj�mhb�)!z���9
g���w������A3�fN��Rꅨ�w��5���$R�/���-��p�(]�TM�-m�Vc���Xp����W$7�*o}�J�����fG&�j��"a�P��{P��xBt�a��4��&+e��>������5l� 8ȁ�F�#��-�]��S��(��Za_m �׷�a��(1�95�E�x%�&�^��uͤ�_ɪ��Y���>�[A����d�i:��5\9)ť����SY�U�_0��b��_z���>��X)�o�܉౒�nā�$7�؞k>ٯ�o���Z�bS���i"��Θ���p�:����ͺ��"+�QC���otW�At�\A,&��D{ᦥ�n�R�W ���_��8ۺ���	�kɣ-*�;|x��Y�h�Ӻ����]�BP�i��	�
�.����^�%oy�4���~[����@G�1,̯ �k4�4@k;���m�a�-�S�j(N����>��ja1���pYD3B!>r���7薪�(�0̥�r�	I,�އ��-�ޚ��u�'����2ڏ�;]��n��F��,�ԼW���"4���AJ �K�P�?�t�4i�v�Yy�xŬ���d��~��};�����-t�i�-��,��O������x�b�J�vv��J�BﹽS�*o���$��JW���l1�.;���䁣]�m~�8��ǂJu�6�Dp�*�ӓ����.X��:۠.�l<�h
�����m��כ�ٛ��V���f�x Kq���V�u��`����{䇮�����-a������'&L���ƣcgS����pKt����]�,��%D�˒`���,�W,�ލ#}.�g�̱�%�F����^y_�f��/�%ع�$~�~:i�Z�֓M�tfs�d]��`��)����O���PB�p%,[w���H@ru�JI17�ȥ�yqΟ^���qܓ��k�쥁�ww���v�'\QŪai��p	ߐ��e�+~�	6c8�C<�(��G�9��Ua=��Ͼ�!%��
���H	N��������*שˢ;�����Oՠ%�_ВK��=��$�#j�~yш��x�]���YE}=Q��R� G�z$]�@`���ZX��G�Jb��&|h���Rԭ�������"�,j�j�����f,A�7���a�N�m�P�M{;G�,����\0�j�pLfD�z��,�J�!�&�����x�5���xx ���f��A7��JPe�.U���e���OŊe�sJ'Ҡ�:�µ�Y~�U瘱�[KǊ�lA`7�%	���!oX���o5������z��6r�H�%���7S��9fz4fq�c�%q0.g<�BF}\���Pp~PLs3�����Zw�Z���Fo 1���v� �>=�!@��SFY�����j�������A:�q�AEh�_��*⩶��f���\A �B_sZg2�:`��������*O�'
;�� ��6GoH<��O���y�0�����Ť��0�]+z�A��Vd�x}�������Q�}ֺ�+��d��-�b{o�ʗPa�:T�QS8�e2��ڐ�4v��5 u����8�#RQ�\�\mtjM��)������ǻ5�̐�:;�X�*�cD�.���ln��� I�c�ܕ�{��z�9�*&�c�'�O����'ϐ�%ƨ������\U�Ի��$D�vU]���%,����l�ѷ����ӷ_U��*���=�v���6{\���Sk̳����/;�NM�K�v+S����z�{W��
;]_�е�h4���#�������۸9�7� 1�:�vd*s�QO��`�;X~�L�� ���s���ʜ3}����<[C�a�ǩ�.�Nnc7��QAA.Xes�K��ҴC�5��MS�J#r��E2O��F+=l=�*G+;���R3��B1?B� ���|��X��~Wj�)�A��т�.��(�]E/q1f�0ٴ�D�*1	�������'Y�ܺ�U�&��{b-�JVos&Ր$���x���-R��]q�D �"?(HŽ�9�w�FeUe��փ?����UQ�W� �S��Uj���б;Ա�l� �,A��Id�Ɉp�RH�~w��fT�hH�g3-��\�hm���S\���BL��2���0^�us?T.�/��-b�T�p H���YS��Kt)k��i�
'!r�T8���2����%���Y�O',�n̔=��E�"��5��&��
� Y�}�mP��7���p~˯Ϥ[�5�g||:��t��E6��h�� U=��к�R6��]4�H��Tz
�U����y�g�IΚ��@�5���Mn*ϡ�Iw�ƽ������J�����������wh�LP7���T� �3�\)�2g|w�f�N�+����]�A��u�Tח�f��8����~;�w��o`�~�p�n�h+�<��:��t��%�TX`��G	��d���4Q�-><ؤml}�#HM�򨯚p����a�� ��4T�DW�H�ભA�C����Nf��3������qI/,�&�6?�F7�Ӌ9�q|Lq��{rlu~��)�KV�d�Z(�����_��+�"Y~o^J�ڿc��pt�Ǵ���2c�#�|sA�FH�AW2ʣz�D�ǯ�ţ�H}��ߐ � ,Գ����(��
 ���~K�t�"���8���,:Do� �6	Dm�ߢ���![��#6�������?��4X�M�|0�@q�c���e�4u���*�9&g���b��}�xr��2<y�e�D��E��>_��V�j<�t�;N�%(-��~<r�X��Iܰ�K�N����� ��#\�V�2�������
�X,`�XM�d���/���`m��X����C;��gD\��ZQ��Ѷw������Ԭ�bƝ�� �ZUGq�?Yf�:�sC\���`Q���ͦ�p���*��Qղʴ�d �6�p�8��#�޿ys�x=��4NZ��Pr�2i�{�ҰD�d�������C��b!�H���95g9Z�D��]�iہ��$��O5��"N
}��hp>7FgݯkLH����w��`s2����:�ąלx}�����SM]9����4��z��fx�VG=���ِS�۰T�t��۔�<ɠ�+Ǐ4�e��pr9��B��j��_m��edM�Pmu-zSu�U�]P#��K
�)�@�ux��$=w���#�6c;a&���0�U���'�yp�m�x����`Ԍ*��r��;3��أ(��ظ���W�p�I����a�z����$O�~�� )�/`��56vb���tB���#*
n��}If�0�SJۥ+��I�D��8�q���7X��K�0'�t�8�"h�fî���Wb�cE'V �st��?�DoJ>]��?��a޹����=db�u(��)g#��Z*�y�NK~�"`�K��<������~����ڀ}s�nG-7�j9���h����+:ٵ2vL�o��W0������"���yB_	^\=��P`�}��O�6
��Pe:��b�R��5u�� u��ӅB��hL��3���>�Aj���W�$>�1?W���ф�����B����xY��A���3� �̌]ٵ'�~P��οR�<��#Gı�Ĉ�����F@f=���G֒{\�C��=]�lFv���AHOB ��kMx���<��lϲg�Re�$��80�͒�
�-���7�XlnZM��:���Ka��M�� '��*�CR8�����\��b5m�Xȁ+g'A�ͬ��j%��)���I �O�UL"Ї׌��<Gk����AmU?=�>�H&�c5L�(���w���.{a�o��a��H '���J�6\}ë/$�߸��hM�r�<��[�e]f7U��u�0��c�ղU���K���;����6j;Vy^)��D,4���yY�= �[D��UjF���x�����t����_6 �ߨ��߀���N�p���HbS�l�t���g�p�Ax��/�R�J�o?�@�X��<�k��W�|ٯj��{�# f� �n�>�z����ǗGv淫S	�Bg�^��8�z�5D�/r���A�$���Ay��w�$����4�Nh&��m��&s���8O&�s����	=�|
�Nd
�R�����1F��BV�oQ�p��r1�l�s��+�T|����x@��`g���)�� ���F>e6��+"Y�wBP��v&c��l�H�����+�f�\9]��q��_i2�TBQ��?O�hRG�jbۯ.tY֨f8<Zɪ�h�0�M	%�����yf���s�Ɖ#���UԼ�t�L ��?B|VFz�H�㐋��.ksG�nΝ�ڂ�V_���^�o�����u�2��KC~<�]��@�;����R\r��k!�4Kk����Ì0�vV�t:~f��6쩷j_���1�5���,I�ᛮ��%�΀B�cE�6 A��\�  �u�;�E|R�"�c#t��t������:,��,,�>�͸afN��[��
���!��r�Z�^��[��K�o_F��6f_�y����*	�6�s�����9���˸�1�]�r���?ω�h��0+E��f����:��,�W���t�#8Ym
=l�����
"�az�o]GOp�,��A�-��:[�K�I�u"V��� Oo���z+v�s6�*��{�GE��l#�^㪍����8(�S��ELX�(V'K�O�eιdT���<�FΤ4�:�M�u��u�E�O��F8�Uj�=�����G1CL$A���:�y=�5n�G�����Vl����3L����LwШH#)@J��A��Gl�` ~��ٗ!o|�!�,U���*ϞC�*���ڞ�w4{\EV>1&V��4[��f2t�hr	��d�9��=SS��R?���z�m	���xJ�+I�Pp��"���&���vC^���̈��g��R�$�m��������{3�_J4a��֦,���m�[�w�+1�I�X�U�+�����&l�y��m���TS�����Ig[����2��A���H=������j(��KNl*o�e������R$n��@!��@Tjc����ה�u|�*�Z��cjL����2Cf�ּ��{���d��:|�?�8����g�fI���ئH͚p�+~o�i?�1�n����@r�>d�˶��F�ڭ�������[CU�F)��B�ˌ��DV�6YjdO�����y!�,K��aj-62�)�i��!M�AJuE�֥+�v�Ԩ�"��h��qT�l̔�-�?0|`b	7=M���DR1�_�R$��#�H+f�h��I�)���jЬ�<Z��w�Y���D�0�lC.]�C��S���4��6��ɺn0Q'Q�+7Y��E��*�0�V����"�O_}glb��n�]DK� �! �/${�@ ���g���럚l��� �z��[���'Mhۯ��3�L)"R�5I B���Zmn4�U,�*�R-���,�4��cj15�X�{uD��n�M�0