��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$��7�4��L+Q���+2�"H�������v�ao4��	�u��=��d=�>�iV�f��l0�Zs��7���~rM��U�`���e����K%�u��ݒ-� rā�SZ )����C.��&0C]�-��[�3�-���+��պݣ�k�J�vo`�A�����f����u�X���v�=�а���]Q�Wۿ�߸�=_Q�X����j>��Zw�K��SvX��ƥ.���#�����Z�0���#7{��\S$��@1I�QX~TQ�E��db����۰� ���>0�%�9�j汈��}��1� ��2���h�G��SeY�a���	'<x�p��k�H`�H�j^y�0�s�78+���ֳ�`�R3dW��_��{p[�?$�s0��#�zS�_��bH
�c�p�IL7]� |����Q�� ��Rr���=��E즕2%�����`�^��l�q-�]�p��jf��Ӽ-f%H���ȳ�>��+���M�71��4_�) 3�46h�rb�J�W� k�h~K0�>P$�_n)���5�r�j��W�J&޴o��$>��6��ŀ�;A~<6P��K�~��f��*I
�Z��}`q���ApC��n���g���3��-�іrO�mF���,�$��@�BI�q�}��Ȥ֐����î�䂧��@������U���vU������ �T#K@f�㯁����|95<@���+�-�)�����K���FI�k���*@�m&���
���ma1[�2�u�I�\�U�yu���o�|��2����;�W�W�}P�K>%5�'�8���׫=����k��,�t�M�0�8]q3���N���GvZ�i�+ C�e
��Ќ�S�v<%���q��e_��
�k�夞��>ZO7E~��5k�TW Aod��eE���G���ɑ-'���?�G$����ќ����8ɸ+ 5ʗ���l�d��,�J�
�^�3b,�����J����#n�zK����z�&��;|�\�^���'e�W�����">�w*<���=�O�V������0g�R��6�c��3Q�<�Y��,k�J���Z�w��Yk����՜@t.G��X(��ї�co�|y���t�g�P�̉�1ؘ.��&��������iqn����bv��Vb��&=�Ě���n��x�0d_a����~ �=�av�u~�ֽz��FBc4��K�峁�9���rdcX�$M�Mb	����L�̷�<�%�G�2�<��ߴ|��9���lk~}�3RY���b���K��!�*�$w?C}5sK�Xx-ȿf@L
��S����)I�Nd����H-������"�e���Y���_Cn��+ViD�;cQ2y��t�c��+~M��	hb�G�w}�ɥ�h����ҟ��p�z�3wA.�w�{9w��_A'�zy�d��5�q�(V��}�s�C�2�;L_�
��:�-:Dp�+`m��;��v��S�P���,n��/}+��V�4�����Dn ��n#!����_4�<
]�����:��u^�t1Ѫ�2�<�zw��4� 3���r�s�LiY�s�#-����`��sD�aqiӧ���8��D�gN�L@'��Q���k�G������v#	��F�ȵ�P�&����f���݊_T'.*�8�)�$���RT(?[�ڇ9kHR��C��F���A���"��P2���5"�ӽ�c�S��@ܬb(�a�
}�{�b/W+�e�4�ܭ̼��s>sBF���.�A|��ꡖ�$Y��=�8�7�Ϙ*�v��|�mU�u��ŅJ�0�I7����1~R�Yhy����:zÖ���l]�GL�c_�8���|5I7�v�yx��:����x�t��m��� z�p1�{��y]���:k��/��1}�

����Q�b$-���+�!�f���IG��e�Қp O�d#Ø����ߪ��u#�:��YI�dp�j�"kM(X �1�f���.�5b���f�9>���#�C������6�!5D�=�Kot�_m֔_��p��0��SUw�������&6\c����._h^�JMS���l2�v���s�`�*�gH�}kv�ل��`LΟ��K
�'���D���ҵ�,��u�R����W���O?"g�aNM��{PBG�T�-P2��=��ģ�����s]����P^�[̃O@׉~ɠ��[�('wfw�_�"N��z���O��V4c<@�ԁ����?�p����{�[�G=<�o)�;�V��E�
�b%�2}~���Z���L�A��C�/��2��[@Xx��(��/ii�pe��.]Qx\�ޱ�� �>�@AD�8'��I�XD5z	�����"���R�q�V��,J��}���4�ĚN��&*c0l[�)�c��"�U|)Z*3I>�(��1!Y7�š�$M`x+��*�
)��8Z�0���2u�?��oJ{5Q�,�����j&}Y�� |o�}w;@���}�2u�if�,�$���HƳe.&��/���Bv�8�{�RY,숋;II��y��>����4f��mrD�e�$R�hBy���[>I1�d�a�?�H4?g�Y=343��2�l?��P�����P�ѱ�
����L2���^�o�*6]�]6�"͝IPsL�j�{���g�	�4È5^T�PFJ�ڠ|P�����1[����2��-p"�z�ՊW����s�A��d	�4|��&�6��F��*rWȯ }��ϴ��:O�R��ASQ�ä���U���-2�>?��c}XX���B�e��25S��5 N���<��q0�˃ͮ4&[˗	��-��PiH>`n) ���U�?^VѶ�MU�9�-چ�n��7�B1��^+-|S�@{֔�ɤ%�����ϒm}}y?���l�bI(ك���r�6����t�P��v��,�Z�@�h����d�,f�c��)�hD���܍�[w�o�ujJ�M_�3
0�
dLq�����<�-���M5&�OxoGi&$������'{��E�+�L��वsY��C���Ct/�f}���{
��@&��mۜ(X$O��K���]oiQI�Y|���m�s��'��"eŗ8�6K���3sh�bd��ӸE��z�f�W�b��e�Ȩ@�G� �z�	����[n�~��>f(�	�����$��m2&���St�d\(�xF�.��!�M�:���^&$�/�F����������Ȼ�T�u﵄�E�TW^1��a�͞����y}F�)H{n+�]�iv<�2�XKǆ��=B�Y�=�j�G�QӦa������a�N^�u0o���Hh����	I�^Pv#���q�Br�O��|��4I���T��rNZ�U`g�/QQR$VE2��3��+Yp��q�a����	Pp�p�6Bz�z�hNS�`��}Lm��x�2����'��m����G��_2ETڼ��=�&/�� �ꚬ��ݠ���n�\�@�d���T�cw^��β����уޓț��'���<S�+dH﵎v]N�'k�p�G�;
�c�I��Ŷ|�Ls(?L�����+Deu���k�^FN������ �P	d\���j����Ȍ�­�&83ܗ`bG�]n~7�޴�6����LJ6o������V��u�5���P@{gt�_Kq�i�y$�\��*���6�>+k3\�)o�g~�=�֭5�M�{�I<L����W�]��f#���7�����uq�E!P���5u���G�x_�KCQ�f��T�?��?�'���,p�K�� �;E���e�d���)�w�"��%�C�Ebw���;�"�wD�f���Ė�\'{2��`��/�+rT81_./������͢�(QmVgZ�� ��ި+��ϘA�����0��c'��[�Bͭ/i��j=:���E} ZW�n����!�V���䮫]�K��W0� ;�{zB3�_�)\
�>��Hb���r]��@p���28D��x��}�_ν�c�Rm-��SY8���ձ��r~��5���ckim��qoϙ�9��6���/~V�ޒ��M��[`��:RlH!.Ԡ'/ؙ��)��8�'����nFK���g�@R�l��aw~�Bm$�Lh���4��++>�j����Pt�kN������p�Y���|���*�� ���� �2��[����Nu�T�����y,۬{&���=ЕEL��	�dLk����������Z��۴3���&ZŠ!�é\38i��fՄ�l���2e9�<��n�R�/��"���$8�Vq��x��n�7X^0���U;��GKW`!��#0poK��U�6%�I"������"�����;�4�}x ��~j�s;��=,"�U����(1|[��(�l��V�tx��|CC;;��-Aߥ�:�a���b�
�Q�T�.�c���{!��\=��R���n��5�G%��X_b,WY�q|aI�nN�FzL��c�D��hI�����[h�z��A\|�iו�h�2�A�0�v�4,xR�r���a-��~��BI�h~9u5�3��|��*�1�ZQ��6��u�m�eЯ!-��0K��;��#Ī�����kܡ�����+!�3�蘿<��~xr�'�%���6�*����I��h1i�<�vb8����LR��c����/D�I;<�0��#[�O�g�qYIz�Kcit�t6�-�(����M�#̣k�M�m(�6�J��F�[dd2b���5��T�����?P:G�,x>@������'�{�f,�#^��M�aV(�˪.auE�d���l���=^h9h>�`�,��(��+�0���P@�����= ��p25#sd�o���:��i�G�ǔ�k�B��f���{�j�I�[��9��N�P�2�g乪��WcQ�o1*B:ER���z�
���1p�b(I�I	N<�%�c��Ch��uXx�3�~ i��BXp8F� EBٖ��SI�ɣ���=R��5��yF0�u�c��J��,���lHGU�.��$1"Ԁ������r=i�%��h��JR������f��D7�
(��Tp�o61^yil�mW�Z��DEI����Ar$���t';��rz���Q)���)�+r5I���sOo�EL�K	���Ř�F�|�t������Z��������[���h0a�2C-+]�vk@�~��)\
p��oI0W�?mɹΡ�d��N�cY��.�M��G	�2�������du�"�e�m��l�\uC�ҙ%�gyۻ�<���HV'�v7��.�C�Ӂ���n�P9C��=�V�OC�}0�5Q�@��%cX!��Ε)��i�mV5V��"T��r��B˩�W��,qN�;I�zAH��L2��D�!�ׯFP��W���\ö�Q� �B���:S^��?��,���dSB�fˈ1=j��È?�T�pM��<�mk
[�H�B����ҏa�h�t�o�%�r���a�i�Ǐ���6}�L4��w?���ECZ��CUQ�E��j��=r��8L���dBF�P�Z$(�Z����]y�K[��в���l�-� ��B突v���;��0��Q�II:�ʢ�����&��PЪa8���|�-�U�}:�+J���,�����I����g�_�����9W�A����o6����,��3��V���"�!ȇa�!�kp?����&�g���s��������L)�3�����Jͼ I"��k�>mq*�) 4իNj�����0�貎��$���nէ�e�;�x|���O�$�*��s\A�9o���C�Z��+��(�J&�)���jر��+�I]jo��kg��<�^��7�
X-���=��P�!&7�PM��cT[�oe%�G-��l��O+�|8i��<�0�z��me���F���xXl�c�)��J_��Ԕ�9dL�:�������,gK�y��R�y�gm�u����� !�B�2m��sE�Ψ:��wD}v`A����+�Ew,IXӥ�č&/��Ԫ�0��fn@�^�{I�[�5�c�N�����cXbė]���΄�G�c�H$OI#�6����@��o^�,)�m�������\l�
ہ�|y%8�p����jS/�j��2��x��g���Z�Bߧ�}�6N�ӀL&�!~���.*�" �z9I�+�i�)`����O!<8W����f�ƍ�Y��8��
F%���؃�ƴ�-�|@�ݭ��>V�M$S���G@VaZA?Nzs�+���cuh�hdd'`�z�L~Rd�a��G��]�c�8�"1�G�B��Y���k�H�Y-������gk�Y���\�@-j��p�9L6��}K���rR ���/�q��ؕ���")��� �連�)����_<9kL��������i����� '�r��e��h.�c�/��� ��?j
H���-(?T��$vS`���`�Es:U�6�ޘ��G�r޽*:�S�8#?���e��y�3{Ȁ*dҷ�ܛ�,
f� 9a}�t���?����x��l���jԦ�ä�K�K��������y��:�7����6��C{�� |�I���?������4�|P:�M8l��p:�xnܧ�]�^��VԼ�~$�9|rے�F�����B�e��erZx��ʚ���t=��q�-=�ǈV=�gy8h6,=t'n
�ڐ7�`�� ��^��V���Pkz8�X���H�&�w�⊬-GcY|����.[��P��f�����M�3oՃ�NV�	��m�;�p�ї!� R���gl���l��W�a%�]5MLf(�Ǯ�Li4K���z��gZ�9w	��릊�<�N�#`j,�!���N
�$)"f*�+e���g�կ{���� ��s"_�S.~-t�+���pDf��W����������E���S�;$v���a̝0�n�nͅ�c�^Hy[��2+ܲ ������Iޛ��K&�2ժ��/�c�D�[��}�_�a�_&G4�|���҈���J�0B������p�*��|P��ſ`��f"�9�GZ��@�]9�6��"i��e�9��y$:��8�2ɨT����Q�4�'����xJ�k�iY�K�$Ӫ=^��$�b����K�e/��-u5u/dM�u'� �֕kUmht�6H�&5@�6l�Wr���Z�V��Ct��p�!�����+]P��փ-����5�
2�����Woz��$}������_
0-ײ�R��;��0��r�LcǖQt�O�B������!�����q���/��QZG!�i�K���e����ȗ!�lM5B��P0��40y󎜩����n#Ц��n�;v�&�Z`�,�is��Y9����S�F9�>kʫ�B�"@�}�T��'��m5�����\w|��L*��
�� ����M%t�q�d�8$2�f�j��=��?%ޯ(N�֫����n��W�������탫��|wޱ��)`�R 38/|J�-�������O֏��T���
��O~.� ڌ�~��9�[%"����N�h�p��Ex��*ܒB�v��9)M�"-DCe��`,�tr�/𐙵>�bl��k)`�ĕ�Bsu�)qcDn����)pG�[ʥG�ʄ+Tm9?D�2��q����)�e�3j|lK㛏�ozm�KB�Z��ao�ŢE;i��W��:���N��Y^�*]�&q����{5�x�r�j�+N><��D�!{�لgb� $�4���b��`��-�&�G����0��{_>~8�D��u�+(6���E���~��ˠ,�D𠨥B�HG��*I���8�6cH�~Gy�=�	&��>�����%�u�nv����g�/����)���t���%�sCQ��RLכ�<}��kFL��	����E��*[����A}�h�=dw�0��������cH�Z/k~Hc�c� 7��m
�`����`�W"n��0�׫7���c����D Q�'�/���h
�SHA���G�"��0��*Kum�}�\Ӡi��4W:se�?��斶Č��%�6���ڶi(h>���f����#r��M3HD�4˱��i<��5ʜ��L�7P	N��v�N�6KSlji����
���</�2Q*�ꩆ4��/�~;�UjhL,f�� w�L�AX&��(&a{�Tx�.C����<������fz!�^�U��u�g#W5,Hi�/�j�8����~�,>�OTg��+��;�Х��E�s%5���v�)����6i�w�<���m�kIڎ�?�����o�#��rᯞ:�
�2��l)B;��hV��x�Vv'
�kkj�dc��q��#q�Ƒ����HN� ������9n�Ήj��ͮ�{������ĝ���^N�++����+e�ǭVZ�7��
��SWG-nW�z�C/r��V2��-oTL3���V$���C=�(R{@{Ͱ���/��#�N:�N "������3(��ԕPc @��Ѧ�����-CU ��"[��@����T�X��,�r$c5�*?��h�r�yg;eg;D��o��V��0,��@�	�����J)���,;7�<su��/'��G�7ۆ<�L�������x�G��iN��,C��Da{�Z���4�.�r^gX��=�g��k��.�:eJy�>ܥr�n��X����|��@�ϡT��9l��F�k�2��GJNh�j�S������r��[S�B!�/m���@[���~����Z��H{+������o6�����z���Z&W8G�|�b�'��90"�뭁$M�W(�u��{�=U&�R�#�q&��*�5���T�U�d� 5Jv?����X󎏊а!�fk.ԋ�AҟER/�h�_t��a�� $Q�Ԛ���G�#�h�E>\�0%*]�������L�Έ�"�L����5~�>��;6�U�UG�6 xT�i�BZ�	��!2�;�1Wqt�v�����C�BH1J��f#��8!�Q4.�v,���f�݂�}siy,l� �!�C>�^sc�/3�"����[�iO8�� D��� �Fr���e���#��73�{e�>��/�Y�G��Xk=L[�̮dv���$��S����}j��[���9�4���h2�}���y\P�K5/J�����-A�n��a�=��]/��W�ѱ)�˕�\4��L}0d���X��B��p��xD1@R�8��I��?@L�(���XL�ǩN�����ֹ~^Ya�8�3Y�+Т{��RNy|A�i�G�a*N�WH�E�`�HX�����?����!#.'�Y�HO�R
�D�*��Y�145�(]��,��+Q/��M�W�>���&�Se�3)�^��@��P�R eQw#ёH��K��D]B��S@l]_�Z���1��jÒoI���ܰ���6;���I��P@��Z���̟�b�^�R-�K3�깮!�弨XȎW�
X�<�=��45C2�54~ڱ�5�B�����S�Hl�ϥ�ܵ�%�dc�W���O�������+�ƀڬ�?j���2�7&0��x���Piq��88���b��|y�6�f�I��2�p�kE�ol������� �1z��ʨ��:��o&�lL�#-^��y�bN���\~�F�(I�T;̈́�jw�s��r��!EW��D�������	P=w��W��-N��4���\���"��%:tC���	~<���*�>��n�PI�G��`�F����%���*{��Wp�`e�������[#;E�ȬD 6��'6�d(�9& �@���1ѷ��$?���F��[?@��"��ZϨ�`%ܷt����"�"�a�ճ$m��2�3���D�;�ÖS˙��4�i�� �qm��F¿��\��9N-�T�f���u����;����G��i=�NVN`-O^h�1��*�q@���~��QI�.sQ�v\��o��h�(m��j�G�E�H)n� �(PluZ�4S���7a��4�(��ʔ��`��{�GDp��6�1��D��
ě`���7�
�r]!�Mk�ϧ�@:�g	�����>��ޫ��=����^�[ъ�t)�����x�^��?�q26��s::����g�w��Y�{Jg�P@�z�b!�i�9����8K��~d�TO'a������ie`�d!6̳�Tb>Y�̱5�X�4�_�[o��T�v�c��g�轩�s�f���#bf�)8�6, |���L$�N��w�1�5=i�
�2$�V�+M���`�kF��C�㉺�ڨE�<�k�����6ޚj���hr�B���� ����θ�B��H����{����;�k�k�6���/(��SXx�l��\�-��0u�(���H���i�k�~OIh"7����)��o$ �,,K��KQw�`�|Qof�� ;��;<3lx��(���PoڗBҠH`*���!��|F�%�U��I��H�S���߾�e��� ��;��AjRO���꬙��c�zE��&w�f0l̻��Q+ɁT��g���L)7VN�gQ��GqH�4A�^��p�����p����2(䤃����:ٲ�9DW���E���@t��uj��+��о����Λ�(fO����Mc#� Aw��$����#ک���:=�^TQȗ�;}F�����=.v�W0=���Ý5�{F.�g��+��� ��Uf��j�H��t����>�N�8m��'y��x m����1�6��7����l�I�7�
M���w���/��\'/�k�nS�y�v�|0�4�����> �jú_��#����:_.�"(V�s��&9TS�fl{����^�Ԁ'f@..�)s��BS�ga�ކ|�h���t�H<p�B�`�$T> դ�_���:?Q��ҡ
Ҏ�U�3�N�t�<KST3Ǝw����>����6�1�{ ����pny�Q�����*��u��i�A�MK�/e�5�����ۡ����)��KǗ]\DLk��v��θa{���t5� W-�EA�
�frq��;�8r���x��dW(o�T�H��_��;FJ_|�HڲV�dƫ�=�KwP��*��iK?��#C� e�t8	�!�����L*��*�����m_�a{x����Ox�8�}�D�dk�8�e ���8n���wЃk"�3/ӧ��7��u��͔O�.`�N�y��#|����W������"a���U�]9ٯD��	��d'�N1��2D�ڡ��zkU�� ��Y�0����QSbU��B,�l$a:��9��'��߈���}��CW���۬��y^B�쥬"�)�ZL�9��5�ASHb���<��>n�g��[-&!f��l9�MǙѾ�<�s�}eg9b����*���+�h9��F.���	��I|o��a�(T��z��ˮ���T�d�A����}\k-�K�&N�L� b���kCՉE�P1�Mڃ˒���vJ�u�V��rMU�}K���;��F�-���H�׌nl�)S@��y&��j������֤���[��v�q��U�|B��� ��x}�3�M�\j�/#s2��`0@�8���p"뛙��B4�+N�V�����i�M�����SN���F6���=�Y��,g#O$	ʹ���f�)rrc>��XJ�W� �V~�´;iۍ�B4S��X%~/���L��d��R4l�"�9[��R��('n1�/��>c-Iq�?�]�*���l��L��TRշ4��O��V�F����NY�;Su�@��V�l �Tm���[���>4��`����<"M_�,a�A��K�+
���̑����`y���T�e]�F���r��0�opZ �W�#'�).Z�|��"I\^�
(��d��DO[kj6�g�5�t��DN�Njr����<!�0"c���"���ެ�y��㢃��ez�"�:��~b������l�.k��9�.Rꋨ�_Il��5��F���E7��)�@� ��|���F��zNr3��!�}�(�S$���Xcx+�n�Gn�%� 2��VM�;�C�`�}�S����������^��u�k%1��E�Xܓ���*Tr�l �������s�T�� Q���u��ޑvIM9>�����ݭl��c�8ي������6@t����b�J&@^��J�~;{;���p]8��܎�U�l# �F�7�~kbw�rv3�H�yi�dI'0