��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� rā�SZ )����C.��&0C]�-��[�3�-���+��պݣ�k�J�vo`�A�����f����u�X���v�=�а���]Q�Wۿ�߸�=_Q�X����j>��Zw�K��SvX��ƥ.���#�����Z�0���#7{��\S$��@1I�QX~TQ�E��db����۰� ���>0�%�9�j汈��}��1� ��2���h�G��SeY�a���	'<x�p��k�H`�H�j^y�0�s�78+���ֳ�`�R3dW��_��{p[�?$�s0��#�zS�_��bH
�c�p�IL7]� |����Q�� ��Rr���=��E즕2%�����`�^��l�q-�]�p��jf��Ӽ-f%H���ȳ�>��+���M�71��4_�) 3�46h�rb�J�W� k�h~K0�>P$�_n)���5�r�j��W�J&޴o��$>��6��ŀ�;A~<6P��K�~��f��*I
�Z��}`q���ApC��n���g���3��-�іrO�mF���,�$��@�BI�q�}��Ȥ֐����î�䂧��@������U���vU������ �T#K@f�㯁����|95<@���+�-�)�����K���FI�k���*@�m&���
���ma1[�2�u�I�\�U�yu���o�|��2����;�W�W�}P�K>%5�'�8���׫=����k��,�t�M�0�8]q3���N���GvZ�i�+ C�e
��Ќ�S�v<%���q��e_��
�k�夞��>ZO7E~��5k�TW Aod��eE���G���ɑ-'���?�G$����ќ����8ɸ+ 5ʗ���l�d��,�J�
�^�3b,�����J����#n�zK����z�&��;|�\�^���'e�W�����">�w*	FO�Δ��v���I�h������l�5����_���a��R�8N��gk+����Ⱳ_�U�ں�H	�#�y���I�o�4��_�-W���qé(�b�n�	�l�w���̃9���[�J�3"6{�Zs�� ����U���]�x���������J�ŪTD)#��d���~I3�LStX��ޯWLR�Z|i>��ה-/��U�B"������K;��tK��������r��6.��psU3Fz�#`�d? U		5l	���{K�.:D���P����r�`{$U�	��l�XJda=�A�����n�pQ��*fw�2����V��������}��:m�>��X+�Τp��I�l�2��PJ:�ݣ|����m�==�̘^1v�'c+��L�3Q��CƩk�@�ι���iHk�\ǛŀQ2U������.�U��w��;}DGP·��g�\�!yZ6��"�ܽ�ZǦA�|�lC[Xi����P:E7�$��~\sU�� X��O��K�bh D�P4����a|7�~�%���!����I;������!D���~L��e�94{i�o�Zχ�d��+��uF�W$��x	���c���`���?M:�C�D��	Z��.Ō�J�y��I�KiW�p����I��7�!�(%\8�)o&����%M�-CtN,�XX���㾩��̯�@�>�A�e�R
 ����S+";r��EwM{o=�����")a�X��J��m�����c%�ˡ��Vn�o�Qt���j�p��g���G=�h�?C�[d��v��!L��_z��C�����t[����L�,��.F��}""}@���3�0��-ie�CJ,�� ۟V��v��3���n��~���B=,��d�m_%NݶR{<�������p�O��
5�#��V�ݹ�(�%a�` �5<ًښ���A��:�ך�r�����3�%�k�R��l�w�'�Y�$���]��?*Gvޗgן6�u��5�{y-��l���|Q��YW����Ee�C�4C�&�ND��e>$�)�p�*�!+y�5Z.��������{/F����++���X �h�5���D'���C>k06Z�^�d5Xs-['�x'V��ɞ�#�'d�Qr-��Ȇ�Qm����p��Q[ߍ.��v��NCJ$F�x@�lՆ�CO�/�w����M�f��xPK:X��`�������̕��6B$U�#ǘ�%�H�
kT�b�:�]��k�v��݂��Ɨ|s��ŞzYR�o�H��*b�e�����D�/��:��T`j�?d�M<��AQt=A:⹙
�ȩ��URAy���x��r)�8�s�#����1)��)}L<�Ӹ�8�ߥ8IA<pEg����a���B�Gw"C��ڠ��Պʮ��q6�����Z�u5���)?�h��$p��Z4� ͏��n�΄`ZQ�[�ëD�$�/�y�P�A�k{*�.��=ڮxq g�c���nd_�g�
���7!��ŝ�����cxqS7j��}�Ŗ�I��`���f��eAA�J@���t>~��~��M��m�jVne�E�Տ��_������k��^�uq]vZp#X�m�R�ۡA|[46��3��2��Q�c"tk3��Ln'�@3�|����m�]Aǟ(�^
�`u�>�Κ�I ɽUG�-�������]Z�nВC�$ڻ�CX�����FL���V9t�xZ-Ç׊˲�㇃��c�2<�:_s���J�E ��>�ܛ$�)���n�)O͚�����-,G�!�!�� D�F]hЎ�DVM"%��F�e�2�e�a̱��#,�`��D�)f[ͧq�V
``�
狅9�" �_g��-��� �F҈�c�6�|gB�>�&�Ŭa���@_�"��" ���;P�	ʻ?��4�ak.#��-'�v/��%����I�Gk0
�}�J���Go��0�/'�IJ��m��T�� ��Z0��н7忰�肿��Ü�lN�H�6��l���$�O�W�r;=�I�k:;���L8�/Toe�]��f�e2�r���i��lda�`h�r�"]�b�==u�[V�?��7e�U2B�FhGBd��N�B�ԀU�&"}���n��PW,��f���G�o��H�����=�K_UT%��'*��33[���Z��@�l�F��_�2]���$��]���;6��$D��m��m�w�uE@�]�YI`����#�V1��x��ds�0�a<���{Q�Cm��P4��ʻ��jR�(��}j�@+l2��HTm/��|QpZ���Mnxh��1��D�HzMÇ@�oq�10��&Q�d�N�,`�#��v�����F���E3A�a����:����U#�����7��l�������4�LE����L��0��o)�=J �HF@��B���#g�?��Ġ�+���9)/Y��1A��s���[�5�p#����z��3Q���E:��*��րo�ˬ�X�W,�ɂ�,]�{��!�92T��pt�6���ִ������ӯ�Pmo;W�m�ubγy7O.Þ��( J�L�F�C8�guB�87�w���*Q�'B�g��b!��>�Qx�n`�ХϔN�Z�P�F=�g�";\��=Ԇ�e���4?4��q����Ũ]Յ�0
)���؍�F��m��k�**��v <��Ӱ��0֜����+�Σ[<��y�[Qt��6Ow���F�k�@ǵ[O��InG�cހve�OԗA�lʑ��%R��~}�K�n���/hCyB��ܰ�Mg�l8�:<���j.�ە�����XCrpW�DEv�(�rS����2F,S�ũ�c)��X'�o����_��o:������H�ѿ��๺'�EP�f��XxP��ii�y�裶�]����-�Ox�!����oNz��q��Ȝ�[}qs�V�hm�I��~�;����/���ם�1ARMA�J�T����ݜQQq�j�b9&�.�+$p���T��܇�I-2����9oq�u�|M���kI����q�01�@׀(D0��/�H���=����6�?���q��EQ#�('Q��� ����P��c˲	��D����O(���У�Lfbݎ-�h�rHl��o0�iB�=���{~��i�PrAll���+�o�i��鱼2q�rI4mp��)��Qs��dD\=4nf�OwW%I~����0&2���[u�?�~R³]x��pxŝ��� ��R��7��䖏��������Ni���N6X�򝡛=ο�K�W��o�H�!r��#��ҷ����c�!L�$�{q�e"`��.H��}�(M�^�I�N��y㩾�$[%Bk�ێ��r��k���^H�:K�wY[^�[q'�O�A�Ђ(�X�_����z�¿�c����)�ql"ԫ?գA�U�He�k�K@F�����d������;,˜�;��?Mـ�}fKk��{Q@m8�s3ip�/\�Q���-=!ݻ�"WQd�S�V��n3��:I�ӥQ�	g�*^w���z�;y�16�w(��j��;yv��t��t˾��m*\��J'~[{�����1�7sY��|��<J��=1� �ڐ�efc����a�����'�%V������&XC�%�v8o�D�v��#?j�����&��l:A��'+�?����L��U��&]��X�$�ZDg`�I�L�D��Ӏ'.�fwI���M��I�GF�aũ��D�ؔ�!�������Z��j��Y2���4�A|k#)�����%��Rƭ�"�Q�+\�U|�`�'���]�RWo�MDaȁ�~�v�I���F�W�ӟ��^�������;ZM3�� 3	·U�R�(��:W�d�&�tn~Dh�� P�U/`���*�"�|-��)o�_u3�GR�՜�Ô%L����YO���ć��!z���}?AMJ�{).���;��~����E��H>�t�PQ"�X���p�J=:7�������Ӧ�u�o���2�-%1��_��H0Sl��3��|��%��G����F�E�Q�USA��ب����%�A���Ͳ��э�%�R��0��P$�� �u&.�'m����t���q�`�VVߎ]r�q_��rgb@V��x��I����3c�ivWatB����_q���M���^���2ډH��+_U�-��^��"]�d\=�>�[��t#r�|87c���R�D-���+�F3���xT��`>j$/���EM� J��s]���}'��4�o��1�'����\��`�>�t	5�eхU�:��ٝ���p��Hq�8�~T]�7־%ȪٲO
<��{��)�w9�S^�y��f��B��nb�=8��,.�s��.�YT��X{N_�k�g�h�n��ר(���v�XJH�k�V1:59�$���o-�*=ydԏ���u���L��K���A�x���JN�T]m�V�%�t �3Sl�|V�L��q�����^�!���^�#	6�rl@�y�K�oy'M��ˬ�~*[Üd*�ޅ���O�����v� k�'��Ί�_*t8��?厌�v��)����l@g>��5��h�n���./�K��S�Ȼ���
����׺�(��]z0�_0�
7`.��p�{�0i�)���/@�7P�T�Ñ�����a�����|"<��8ݨ^�6�hl��N��������z�	t�='�s7I`�VKMk�rNN�L���O�.v��Pt�T5��bպti��¦�K��}���g4���S������!�?�aJ�d�;������<4��+Կ>Շ!��v��WX��L. ��l������-p�X3��ig���z^
���K��`������bc&݋U%��-8�Ǿ#?	�2��NهKw�� D���g�ab�������"o9���6� ��&U��N��u�>3���3A�jP����.��mU��2�Z�
Vǂ,F�ڴVH�D8�&��L��ԋ��9+{k�`0J���PtVr����_�n�!�YEeD�9�R|Ά�1Ňx�¬��-�a���4��0����|ם|FulSaվ�8��bOsD�pϮ���	2Z�_���`��v��Hw�:�͔�С6qQC�o�?Õ����Jʜ��F�G
eZ� �3�yي��HW��n�ǅ���� x�)Lj��a���vF��i�̻���Xm�z����ދ֏��z�u���ITI���z�V��~,M99�p��Ӓ�LQ���'�N������ly|�.�3��mf10�ѻ�d������s1?A�NxC�#����@�.�j7E:��SRX|�`�K�B��ךW[�2
�3��>]���|-
��/n��әL��%ܢ��|s�k�t��L� 9,j����1&S�SNB��oZ�MB�W�Y�eX�%tb��:n��`\S�H�n�K��GE�8�޵��er�ԙWa�2��~x� 
�ݓ�����(�Yv������8��}�I��'�n�J�|R_�E�$
f��1�Y5ܧ+r�د -�;T�ïO��n�H����rvآ��UnF�V1�^�N���z���6����T�Pc&vk�fb���Bb�3��T^-=�1p�CS�����y���U2�pF4W:|��i��3E�0��]߆�������M���OoA����'���5(����+&MP�4,#���au�f�!�%P�A�k��������c�H}��6�ŉ���F֒�c��T���#+���٘�`��\Kz8]�0v,�@3��Ӳ���u��?腚a���o-b<h�z-�Arq��L�ua���D�-��	]W�:��e����`.R�	�+�X��*b�c�3k�&�2Q�#�2-ˀL�Pᙺ�=��8��f��@�H�[i9�~�Q=[�m���a���������P���T )��s��U%����E����ڛ�����F-.1r���L`�^�u�$8H�=�DFP��	�xa�䣫5��v�s�JɅj�jၬ���#^�_�c{VJ�;t�~(OM\
TX^�;[�C*�hU������$j#��#Z��P$	Sw7��r+�/r-g�y�Q�4���h�n(��qy����hZ�.��bC/Qx9�5lTnѮ+&�wS�`XN���Az�Bk���Q>Sƛ�t���.'�& ���lt3I��PU�=D���`�{�����9���SE^��+m�n	E�A&�E�[�8aiZ��+�<p��������D�ꔮu����ڮFKm$GEtW�k2U��-�m5{��64��f�o!�;w���о�1v�ȋNNH(�3�*�3���O@�_q"���6�M6������)�]��7?sc����(�'�Қ�{������|�q���4	�,U.��;�CTU�T́�3#�\:׭��r+��fD�GBu�(_��]�{���7�b���l81�@��b�����,-)�h\U�B&�>��C(��"O��P��2g�Os���@)�>Ex��T�]��bkn~E��h��b
�ަ\hR�~g��d�C�<�7��]}��Ko �_N��H��kǂ1��]� D~3��z.���x��ORf���aB�J8�4��0��=��<??^)i����dԴ)��r0������-Ta��He	�J�`��sXXi�͸!=X�1{���s��0hO�k1Bc.���*k���E&�꩸�� E���+�35��k��dL0�*޷�șQ/���y�c��(d���v�΀t@2��� ��<����/?�/�	���)��:�ְ5/gE�V$��I�������Ǳ�(�a"�X4�-�}�R�oU��tLv�G�X_?z��&~e:�l����ٓ����C�Go����si�
����5JPE�[��[��{ ���}�^���P���w�>�S����M��{�c�(�g`І4���n��F��:�qdAn���(疷8ُJ�w�9ʀ)'4�e��������i�J��R������0O�� 3�NX�e���M߻��0`���
������c}fX����dy�:�Zv�
��D�l���x�)���0U����P���]FbEN3��lL���Fq�]�����g�@�v���>y|��G�v+�O�G�9��Ek�������VaĄ�H挾�-S�ss �
n��f��=�7�C.7�Ω�:��F��f�Ƒ���(���lDey|����Th;h�@��ѕ��6�,۪���w8n��e�7�
���U�8��$l�^|H��Ϙr���e�iȝUe��,�M����v������CP.�s�fu��]Qg�u�	"(Z������_Q���Ew*�jǹ�ߚX��~�s7��Ka�S���A}��?l�`B�3�q,�}�����Y����n*�}Ȗ���z�n�I�+@�}z�RTr�3Hd��ABʕdt�H�g��g����nf`��B#ݺ��-*�\�E�?����x��[�h�8�,/�#���G���R�Ƹ^N�5�a�֞�m�9�⡣i/�Y��^�C��J8�(V��>�T����0�͵kS����zh���/#��4CLx��|�f*7�#E�B2L���|�+�BA�����-FX:&o��� ],�ʓ^Y)I^�����c@ `����9���M�ԂU4�@�l�v�{�&��`A�6��S7eD]��t�jx4i�|!7�~㒐��>}߀�����j�.�7`e@.�.�2���8�b�SɃy��{���I�/���{�I��|�$����U*A���f��9����o(���5
�fS�������LQ:��䜠ҜrV��m��x8�L+��(�?]A� }����А�`�����}��F��2
�x7�(fN��S�����~���ä�s�N��Mz&E��*�D�M��ߦ���Z����	G��N������k@O/!6A`��: 5X֟Δ��S�Q����@3���oؽv�J�Fjő ��u-��ߨ$_FrM��2�͠1h�p�½iGX�[��zsJ��wH��r.�R ���#�KO��!�� l�?=����B\�.-�ɵe�O��'�9il��0���C[w?RE_�d��3�K]qK�ɮC+Wu_����_`{�8����;#����i;&�F��� ��Ը2�c��3��7G<�#_6�4�7a�b��
L�R|c������4�3��9M�M��R	3�U�A�͒튕��d+v��'���r\R��ГWV$	�.Ô���\�-W�eϣ�����v�h���%W�,���������Ѩ����G�h�&iG�h�A;W�'/P�PP��ZCC[6��M��V��h1��?p��2�� -%�=ʻȅ�!}y���ʂɀ�+���0�:OB�z��\呂ll��fٟg�_����E��_-Hڦ77ӓ<�cM;p��	B�՚7:h)����0<TyH�	�=����3���/
��{:��T1"����H�YMJat2EL5���n)Y�_�I�`��h���y���.^�6�HD���Ǟ�W�ch�r�'?������Q �gc�K��cp���gXW$h�Q2����P���`P���KV��!���"m��y��L�>���5yz΢�ō�N���N:u��ѪH�Q�pwB�J6�bt3x���˶TW�q#��A�� l���?����_�ª"4l��Z��ۃX%7�>&����<��T��z���oJr歰
���9��;3�e����"M���z�J"&1M��1tiަ8$�?�+%I�����Xk넌ƽK�V*mqd��el�s�eJ��Ck� t�q������=��##�|�XïҨYR�BDN�8b��Q3;jNb��O����<Rw�6��6�����(хd�ݻ�{��Z֚(%E#|��>А��i�f����ޭ�.�W�ǁ>wY�@�R��vN�l:H�^���"n�V�?$�s`��f����VwȆ��×s3$���Ժ�fG�|
�������si@K����
ew�-���r�@M���a�:j��@�[5�y�V� Ws[G�V��GR�V ^?�F�5�f�T����"�Ծ����f7r]O=���_� 4zR(�]�������YbD$��'�Í8�TC�-�� &J�RB���"h#'tǶ�Q���\�ET�=��+�QjP~~����%���]U%�ՖJ��
�A��OĚWU�Ic��gG�3��eA�����(�͢ߒm���;F�ƺ�M�󍠝�M��ɗ�0��!���E�ު.�?&�I���5?;Q
�w��l�b"*{�aP���6ݯ�F��]��p��{�i.��O5����Qt,�"U����S��x�u0�づ�.�Ƽ�5��˺���{� ��� y͕s�~�e��ǈo��ّ��Oy:c;9!�I����$6Եn�գ�^�ID>�״�<�2K��xVdh|�Z) ByB�}�۳�������C���X��6�R�~�����&���L�wZơ�Q���%�nx�Ԕ�L��h��8��y]����J�c���=�?�b� l�$D�p+�w�'��V6ǎ�LT�%��T׽����j�aPV>�ʹ�A���� �$=��O�Q։mz�эQ{��i�4t�|��n�y$��/AVs�ƿ���kW��9����\�Z�D�WJ�OR��R'q��9�^�dK��%:����G���z��>��ل�`t�{�/8\��,n�������olW-qn���z���ӯ\վ�0�`v���Xٯ��';X�&�3�6B�nj�x��-��T\N_iȧ�Cm��A�.�����e4�������-�f�
#x;���MbF卲P ;������'ȌyzP�i��1Y{��L�q�ݮ
�]�kS�!\yO;�v�I
�fH�*��ç8:FX&�f�(|���ɻ�吴���R�@�J�k;���f��+2�C4��x�3s]U��a�=�B2g5\=X���n����i�Ц��6��팠��$��a�=�
���k��u��Pt�L�y;cћF��Sl����j���=��т�_��~g��w��L>��%Z��=�/_��\���w@h ��?n�A�?���ň�Q��7�ף��+>�'\b
��k真� `��z��2P�3��=(��2p򽭿I ���HĆ��Ĥ�ޟt�?��7��s��ר�����l��^�	���V5�X��������� ��by�R×�B-K'�݁���i���<�*�c>[�}��۳�C-��4�����h��HX\��=�z��t�CS�?��I뮴��át��!�w`���I�8�J�'��3�őЈ`��Z���vf�|��q,t����E������o'P�?pc�:�k[ګ'qPK���\J��6N{���D�D٫�t��T�H��ԃX|&&���e^���)=���K1��$xr����Py0����!
o��Ĺ�5��@��EG�2�bʨ�]6Ngc8�2��x{�^�4pM���K@��=^@vTg��q-u�2��^���
io����l�'������O߰���n��N�@�Am�Ub���eۥ�M����6˾���k�+)�L�MdX�H�5͜tiLE�|-(�\���}!��M����3�٠��w;jVW����u��=����PƔGy�ݳ���A��w��Jrׁ�����g�uC����j�\�=�"V�3�o<�h/�Z�s�r)��56�-b���k���J;C��5'��Qq��K�	�K�� ~��,��
���G�QjV+��z�4�X��#�"��C���
��G�5�A�ʊ+ͥ�	�⹻�#RVv���}��r��MF���_2�x��_WYb*.׶�Ĭ�jٌ��af����Ƭ����ƌ�-L�<.T�S�(���*��1�N�c�ź�e�p�������x2�׍�� ���V�(�Ze����@��!����I�Mي'z� j���~���#��;��E���	�h���}s�2�▎ۮ����OϾ������Íx$�t�)�]���#5����&����Kg4�Y!+6H�z�Ot���&f@��Lq�x�Dэ=�wN7��~1\4�4�_�Ǘ.m\{	ҕ����uf���n޼�X�8ɚ��~�9/�,��$F���g�L����v�qb�3Zk�b��"���ƺ567N�����Q��THԄ����Im�#�,�G�-{�U�ܛ��9c9��]�h4{t��-:�}.������<.e�5u�8�-lFU1���,���2�7X����4▨i��G�/)��a�Z�O)0��᳔)�)=��P�P ��<yu@k��e����|l�YZ��2tg���B��#Ϳp���܌����hg�Z2�oN��)"fh
-���_T�͉�K.�� i`]""�Ŭ.�UC�Ly�ب��":ݢ�0�t3�DqԽ�C�U~p�%H�Cd{�ᨥ�`F�������C}�W���/�=q�L�A�%i�&s�k!C��Z��=�Zq�4��.U;ᗥF�Wu+��E�Q=�:0��R
��h��QV�m��+�!E�)��d%�r|&�/�)JV��
��	3O[\�tkɥm3�W��m�l������`�ȣ[�{�w጗��N�jF��H�l]duDc��M�M|վ�o$q�"P�{ݝ���soZF���O8va��-\���F��f_���P)�@�����{ó��5bn�ڡ����APq~�p��r���eX��X�ZW���(}���ٍڮ{�G�23�c��|,�QC?
]u���W�y�����}"�p�޾��@�D� �O菶p�R�Jd'���?��l��[��#�Ťކ'v�&-T BbZFlt���.9�+G5���k4�FDH������"�"�DF�G"��{ʾԉ�K�$r���xZ�F�#������Vi8�������-�o8M��v�ec�\��e�waz�T�>�  bc^��(Y�|;J9w�;���6�P�����0�:�Ƙ����^����k�(Ȇ"�76��ͶH���- �� �k�+G�W����m`��x�O�B�5gyRXI�,��2��w3�-��p��%m�
��o���Ư�2�����$��@Yd4e�j^���Qr}�.P=O�#�H����A�Ē�h�*�^j��ovK��?|?
P����B�#�\�/9��	��̈�����̼7i;ҡ\q��r��T���O�0�f$zh�:�Y�/5�`�Vu��#��Ҟc>�{�]"��%I�2�V}�����I�&
����k��X�pb&�`�CG@��_�Ĵd7-�8t�,�f�[|������5�*���wi�SJ���ϫ�)��C��^�5������{	��y�L���Y��3#t:��Q��~u'���ל}֬���"��1Ǭ�h9&��:�
�=��5�ؔr]��ŋ��;�K�� @>�qwj�����r8��>*f�Cʳ���i����, ,}z-Z�(��C#���!a����8���:VE)f"ݔWźV��ڶ�T��D��kץ`�[N1�JRب}R�ۆ�{+�z\ N���Y�@��j��}�Q��� �I�v��O���V`7�b��I��g�h�	!ys6�L5�1��*s)��eQ!�l����������������5�?g���FB��p�ٴ�3��WyZÌ�\%ɛ�*���\���ϝ"�.��]�p���LCb�&˺S��v �s�w= *6�L�Hn<��Bb���0�b	:B�EU;БE�0ߔ���X{�3����I3�XeG�U� O���������P�� 5pꯇpᑶoYX%���������R9�>����nR���߰�,��x&X{���i������XUJ�ׄRK1�O����e���?F���9ƿ��*��XGR��w�P�f�V�~��t��z#��0�	�Dm�8ֿߌ�p�-�Jb����$`�����TO�X
�Ĵ�Pf:D�0ߍ��(�]Q�v��n�݄L�0rJ���AR����K��eY��]�5�_�������E3��d%tc�}�2���*q�%s�5s�%X�ŗ?�C��G�ˠB�$�a^�Ƙ.��o������c˅��!���ϗ�3�?�J5���,��εȬڥ����HM\����412���"��u$�tH���}��4'����D������O�/'y*C"��9�L���T��px%o��<�~������I=K\O�8r��I2������3T��wd��3�@�*a��'
�9Qg$��fap�1c��98��8�����,���&n6��nǫ*�F5�u}a�:���Y�G�<l:0��������D���β�vJ|Ԅ(yXU����Dr��A!D���x���������0:\��瞻\H>���Cz�Wq��)^f�_U��������w)i�{�����Q&!�W9}�
7U;�]Q�3�,|�y�"y6���l�+��g��I�����"~7vJ�<kl6�@mƼC/�e{Q��yv�׬:U�QF��P���Đ��%�O�XˉOZ����C�0Z.[��1%��*d��Y}�jL~�b�cD�md��X�b�,s&���)m�S%�%߳�U�)�:�d�������<��}�#'9�0��:�!$.��n]�t⧂X���g���\F���g��D���T�"x�g�qtr8	A62�Թ'I�U�v���;��+v�^���ָD��no�@Ҹ4�oS����ݴ�]m͉d,���r�Zk�������6����膀����nQ��/k{p��3�q7A�t���Խ*"��,Eg��W�1��f�o�j6�k+W �Y��{>��x?Jׄ9��mD{%��9��i��B=#���\�c-��6���"�Z�O�x�L��F��5?��3��y��%��?���ڨ�x\ͽ�k����i��?~�j?-�;�	IHU�IZg0����A�(A������Ab����#^(	��n��?�f+k��:�*�&�x��H��O��䒪A�Y����5D	+gJ�D�N_��V�t)|�C�t�w���yT�:����>�y�aq�i�ꒄ"C�m7��3d7#H6T�@���}�Dʦ3�ſ>kHf����Gu�_{�(�<�X��T�9(���ޓ���1��Ck״���{�_�KvU��KJl�u-��s��H6{�)��9�d���xwx���u�����z���.bu ���,Mh�%��������\�Ά}�k��d	6�z�X�x�Ve[�]�SoN�����V��:�]�Z�5��x;����O���ȖH�x�i�r:~��T��~.8�~]��F\���ۉB\���IRrhşAM� �C��y��	[��胀z�Q��B	����k/�����c���E��ɞ�qG<���E:�\�(�z��2�>ro�
�k=���މ�0,��z8������uE�´kL���Y�GH����@����얝!��&��)@�}��z�׏��,��;����%�U��*�Z]�%����#���ݖ�-Д���/�1��ڠ!�]$u�<�C��W%�`�R���f�9g+daE�`�i�ic�_�f��3������pl-�Q�n-��WZ^\!v.�荎�G�~�<�tGF��:vh��
R�|g��*�Q����M�򇔂t<�;��0��L|ѣ�h���K�\%���=����V׉��M#M�wЀh��-������f��Q�l�s�#P\m�ڀ�疱*b+��vjC������Cߵ�QV��2c�G?����ѿP3:e"�smٳ�pa��u#�۳��ĭҌ{��W�Ǐ4�뫂v!���>�).�^c�B���� t�,7L���"8�@���[��K䖅��9<�#�<��,	��8I¡�5|Ɔ ���}�Ġ+�߇ӿ�U�Xs���NYnP�r�l��D_uS l%b���[�Ԁ$n�S|��H����u�;�X�%�5B�Ҳ�0g�>���I��q�0�˪wɓ��XqJ�(0���sn.,�4��,��[|.@��Ӯ���<d��,1C�qh�e�t+6Ds˗�3��+��v�mL.�}dw\�&8h8l[d:k� M#P娠7Ƞ�w�8F\9���F7��MhV����	�IǦ�����z)rNc�H���Fk�ܼϱ��Z��+x�k�J^�}�⨦�Xh5���Ǟ��X�|,Wі�(�e�k~���B���h���B�ɯ�Ȱ�d;BH����	��g0ʡ�kT����E!��8G�/6v�ӳ��d��F���8ߞ��}�R�p��՚2�(�,�'nG݋[	V�����C�����2Q3+M��QXg�ޡ��UM1�Z�P�e�y�5�3|0�D��D�	��<Y��`��5L��w;�k��
"�*��A45�8��@�[�l~D^u�6E�u2��'�
��XDӿ�#~KH9�&/T�ã�Y*8#��[� �����"r��Y�?}�D���]�����dї^�g�A���8�C�P/� N���F��q��Mxl^������=�����쥙��DQ��hG���*�)@6�%Ҹ��Y��h����x�]Y��W*���d~�=�8k`����‘��d{?"h;�i�b���9m#P.~��ԅ3�4����t�#�|:0wa��M*p)���0ƾK�	�k��\H#��r�Y�d� /�#�.�*�T4�J�`�S�$L�<[�;j�J�/�M�M�A��]m㘘{Q��I������`˳��-ȱHF5`q��B�fU�G�tvXy��3��ZN�#����(у��0��-D�d�N���̞$�c#OP5*��O���GؚN�C���Geո�Ҡ����}�����.f'M[��Q��h��(@o�(X�\��;����Uw���Pk��k���)e��DQ���������x:l���P"��-����S:3NO�dz�����yJ��K�a��ő�S6 ��s0�ݼg�b
O�+Ͳ������t$T�V�Y4h�雚d����r�͚���&ұ�W�F9�Ź"8%��<^��m-ʌ��^�7\Z�b|�t�_�t��q!�l�l��k�S)KjH*���~�N��`{=�d�4g��?���ld���g@�(>���m�τC����� t���C̊�w��71���ow���YN2uҫ�y���N^�(pV��6wb��Ȍ��e�jr(HRId*����>��BѴ��!��F{������V��� ��x�`��ڨ�QF�Y0�I����dM�C��NAk�1ʤ�HQ�T]�Q~K��e롕��<����B�7K�Ar�Kn"�[��x2{}�.W��'�M)�wi-����u*�R�L�p�T�k�N�����y��@ܫ��R�@0��ZD�Ύ��p��@ӫ�L�6I��y���/�	,e9���Ҽ�"58r��`���B��� CGE!���_1�p��*�d��rK���<�����6�ވ��+���0?s^�2Ȑ��v����<�5�`�7o��~�~-\]���ǖܿ�҃()�\��=_b���������?��ȇ�����D�
c����7}������t�&d��&¨/&�����Y��/G���V�'����rs�U����瞘�\�X�]l��1L lS�*����l���Ħ�6Z��|�`g��;���
w�&����t�$��[[�|�X��9.�h��nAk���0����Th�D��
�o�Wڽ����y�M���Ag�.���h����a��H�%6����\"$s#y)�p��h�#q泆��]�[���=����@K��d;%���u`S���<TXC��^�{2(����Yc���zfav�kK�(!�R�[���������1sLa�B�n��A'�5��D�;�XQ�Яi9a�Ȥ�S:ܯ`�.=D��«Ft����ZHP!��+����M��ANy��*CI�d��i���<���V����NQ;��PZ��m�H}�Ly>�����5�5�K�����=�����o�2��9��zA�I dܣ	��
Q���m�P�~ǯexft#�{b ��F6���h��T��/��ts�x8�x��������~��Dq)���i"� �ju.̉�9t��,����C�N�Ӻ�-�!^�����P~��y�r]C��ˡ1n�����R�	,��S�0ꌎ��rw�����uT�S��4[2��e��SƏ�S�����k��_"D�ڮ�{��RHAq�Ї�*z<>c����L��ѿ���
��*��W�6UȀO$���#���c:�� ���%���@F%�[��z����#�O��^�_x��D��X$��!kK��4U�|?0�"�Pw���=�� ���Lo9��M?�k��L�w��A���&�c��Jr�sZ�������L�|J<1��>t�o{�`Ǻh��[$�o5TdH�f��5�7���n' �Oa/�{�e��D�U�=�
+�o�0ӕ�s�N�涣(���S�;���f	6<�-��;_��-�ӂP�9e�28��оm�+@O���3��p��R��=�D%oR�/��g��T�7YKU���/��pT�����q�}J8��J���r�*��G�Z���q���S��G���F�8`�:�,h�a>_B��]*=A�j�9|�*ܵ���A>�iC&I�
r�����C|ICA�e�������N���T��@� +�rl� R�Z��>Z:O��ʈ�4z9w�Q�_���`�@�_�B���H�oL�ИU�pC �L���ae�i����
�#��%�n��79%�$X�ח��6��]:�cضwՑ�49a��'HH2��.��զ��5�aV��ȑU���zo���O��rķ;�#����.R{��\�f��_H���2��p�S�3�5���b��RQZV*F�?��|��b
���A��v���sC�@��Y��D}?�`��.ېT,@Pq��S��l߂�&�P,!�⺕���1G�#47�*N!��Q��[4�³�s����I�/P��D�kO�ҡ�����{C������"�[���WeĪ��-�9Jͨ��C>���N�R-���-���TB���.��Ra������wv��)����tګ~�bA����,�"H�b�`�c�������� �2�KQB��yƘ�Ԏ�ܥ������L��q�rg:#��<���űg�����5r��Ğ�7S�����K�������u��K����S,˴Pz�k�q��!��^�!��n��q�t&����z�?�����.(�͒{죯�����1�h"q�NάDM*�v�QyZЃ�>
�|:�9SD����x�ߘ�������Ӈ��za27��y�6�DE3~,�_ �4�5�����6�P�{-}�N��S\N(~�����]s����Z|�#7j��
�w�������w��*%�e&u��Ԍč���cG$�|�^j��2?��%y�ʗ�VO�D�<p�Ҵ�?@���[	 ��ď�żɅ���_�7��=�'��OIL����3L��f7��:���䯐*�)���z���kx�P'� ���g�4sY�tQ�v�/�bwH������.�����E�J���dմ�:�
�����@��m�_��B'�[��6�f��HD���3?'��˔�h���n~.E����]��\�)7���zk�����&G}Y��*���&�ɍ�M�Rt{������8���҃7��{Y[0j%��T]_��z,
ڡ뿀��P��wo�.<E�v�����,�BV7_`Xzxe�l�&)�V���yp���?�������U�R�]͚+9{�I M�aV\�4�?	����38{WL+~��#��Z�&�,Mqx��{j��
��H�cq�g[#a���)A;)��[��"���� ubUX�QRV�m]sOY9�E�(�d�oK4��DKGL��F�ѹ{�CY�
��l+��D�q�z�S2P������b��)�r� �
�iL�����T(ELU}����ssn}W!�2wţ������W�?pb�h��+iu]�U\��B��hpt.��E� ����
'P�swjSc�\���9f�jP�>��g��{�$��E�;N��߄�iW���1*���S�9(�[Ho�u^�-�E^?�#Yp��{v[���M����j��ȿ���ǫ0�;y}Q8���hI��gن��U�Q�������jAC9�}���������"y�M�k��&=���ӥF�,2�a����R{h��h�lC$��bff�"?L��f^�z�L��ep�&��&�uG�|y4zߗ��0k �5�K�N^�*6�- ?ϋ�D�R`b���e�b�P�����^��ז����bjF:��i��0~��+S�}����?������mo��p�b��y�|bQ�[{bw�	�/�<N��{k2��)=�8I>t����-ۖ���bgĆ*i^R�k�;>B��:��İ34G岏�&2�ݱ�u@˯-����E.��3����XK���.j��CaP�h��y�\널C�Ϣcx�JN��8��f�3��QZ�#Z��ȣ�+Czo~o{�AS�U*�^s��u�{Q��%<;�!=�.�o���2�]L6K��`j�N!:Ib�[+�;�SJ|�<�^N�!ry����Dp̏�$�
"�5��Y�?J����@��J�E��
�|�
T�:\�i�h�	�b����ғL6@^��D��O��5������1A(�_}�S�$`���=`�,�'��J�|���43�i���Ƒۛ|���LNѱ{A�cSxk����l�3��AY�B�>\��=��|N�E�����9x)R�� ��f��og��8��"�`�%�E-+�z��8� ���=wp����GOG��`礶H�G���\���V��zk��`E	��e\�ϸQ=(��`{�9̑�V�<:�D�n���L8.|n#z���6�$v���- }{�G�;�!@X^ؓ6^��KՀ�-!�}ŶsN�+ �Tu����%B#�m��9^~����U�1rذ��37l�������z�Н���79S������tj�l�z��>%K�6{�"�dN��%�foIE�$K���U�'�Z	9y3���3VYz�|�c^�!.7��*gtl��Vh�.M�'�3��j�{KK�wb��(	y�d���wp�8��3�i����e�/�4{�k�A��Ź�͠Ɵlr^j)��@��v�.�[ߏ3P�Z�w�4"���V�N�Z��R�JD�k��=U�Jǡ�BpucD�ʓ����3a)��~�k����d͕`%�g8E�%�Gk�?�5)s��k�` ���}[7g���pr%�(�ҥ��a�y��$�~˚)R<�ɫ�F%��6�r�ְ�}�����QeN�.�$��?��� �;=�k��u��浰���,
tc���]�Z���ʳѩx}�F�g!3�h]<5����*t��n�� ����o�v1}��)�n$�X��7�c���e�rŰ컞m.�̎_w)��K��
�%T,��Pv�Ѩ���{7`���u7��~:�+@3���)��ь1o�� a�k=l̛��:o�-��5��ɺU�'ׄ *xp
NUb�[�����r�2��L�OP�i����y%����[�5H��AQYϤ�C�����h.'�Q@�%�t�Ad!7��P֟��d����{���K�N��וşp�Fn1F�v�*�e�);�U���X�R�V9�M*�?cybxqd�~��?;��:\^�e����6���x���I��d��>�ȭ;q�f�ԫ'Y�V�=��F��_~�3X�d���.�U�b��3ࡀgÂj��0�|N㝗�o�f��f���!����b�D5�{Qn���wJ`�&+��Ɓ���@�*Q5޹keI�)F�����t����*���A!��E*��/�6Q?�� �{=Yο�����ɘYyQ�Y�?�定ʇ��	فLJ�՛Z��7P�&�4KZ4�"�����.�e�O�y��bX0�Kq���8d�blSKnڙ�^ʳ�W��V��8�;� B�LXQ�#�kn_��F�X�����t�7�	6%]�3N�WI�}��u���[����pz��2)�;M>g	�#��nyȠ�S�I�Dy�_W:�q���I�,�s��*�B��TA������ ���Ӏ����D^I��Io���G�R/��X�Q�Q�VTO��v~�*�pv�'�m���m���)��WFf��6��d9�"\��'=�_yt/y�%�0��)O�J�����E9�u�Nc��(� C��ᢊ�6�[A'ϭ������+