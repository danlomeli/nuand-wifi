��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� rā�SZ )����C.��&0C]�-��[�3�-���+��պݣ�k�J�vo`�A�����f����u�X���v�=�а���]Q�Wۿ�߸�=_Q�X����j>��Zw�K��SvX��ƥ.���#�����Z�0���#7{��\S$��@1I�QX~TQ�E��db����۰� ���>0�%�9�j汈��}��1� ��2���h�G��SeY�a���	'<x�p��k�H`�H�j^y�0�s�78+���ֳ�`�R3dW��_��{p[�?$�s0��#�zS�_��bH
�c�p�IL7]� |����Q�� ��Rr���=��E즕2%�����`�^��l�q-�]�p��jf��Ӽ-f%H���ȳ�>��+���M�71��4_�) 3�46h�rb�J�W� k�h~K0�>P$�_n)���5�r�j��W�J&޴o��$>��6��ŀ�;A~<6P��K�~��f��*I
�Z��}`q���ApC��n���g���3��-�іrO�mF���,�$��@�BI�q�}��Ȥ֐����î�䂧��@������U���vU������ �T#K@f�㯁����|95<@���+�-�)�����K���FI�k���*@�m&���
���ma1[�2�u�I�\�U�yu���o�|��2����;�W�W�}P�K>%5�'�8���׫=����k��,�t�M�0�8]q3���N���GvZ�#z�HM���f5�����;�q��Pj����H�L�}��T7���z@�o	%�PFmy�lc�
)�8yIf�o���Z�"4��r���o�6˦��)��"�~���6��}�pY���]��
��K,�	���1D�̹�@��$���(_kk<| &���x,�u��Sm��Fģ	U��U9�k-��c�KU ��1$k�):h�����!�Έ>�l�B2A�V쉀�#� o�Aڐu�Q�%`��ܸ��cb.�����E��&�Ѯbz-V*�E���bnjۜb>W���z�<\UlA"���i��J��Xj݊���	p��k��1O:�$w%�C�\��H��U���Z�W��k�B�E��d��/���|�0�=o�g����/Z^����X@�N �Y*E�M��j��Ʒ�G��V��$��Qhw-J���,�B�����>�n�N9+���̍�)ТP��yw�~2�]�4�E�,��$&�_�������%�#P� M����PA��[�Z]�ϒ=!�ܠ��T�X�`2s��gq�D���&��%�?�Gy���4E��[4�͹��*�r�S�Q�����!P<�g����j�m2W|���i�:�?���_7��[�@k��v��I�������,��u�T�䷏Cë(��5<-�����8J���R�[{{l�Ijt�d�	0�:�K���}�� ��@W���D���&�b�kݿQ<
�d�dl�\aJ�n��En�V���pT���u!=��$�Z�
���Ѭ�!���w�*� ���NثE�_ *X��F�A
^�7��u ��*r�ܜK	���7�,+�iպ��z��<�7��x�j�ԡ��ܿ�bx2w-�lvDd�T���$:�k��l��Mr �n诗�Tcpb������/��h&�=��|�B"����Yb�=���t-�B��[K߹�zKVX�ʳ���_N��hF�Z�3 �<�~[0��s�ـ�`��=�sZc�B�<Q�"K�;<�G��grN�4�,U���3:&��w���"�p�`��u��� .<����h=���N`��G�e_c�\T,����2L��lއ+U���� |��!1K�߾������6��]�C3^�m/^��q\ �;>s�p}׀,��3�w)��
��q�7M6���W~ �L ��J��R&���@��}P����^m�l��@�	�;>FQb��c�N�>Y���]�� _�����;��YZ�K�.�F��*��΢F�I�n��x��xK��1���g���F�J�����8�:-e��O���΋�H�K�g)(YLP���̌v�)� ���9�l!�t���-��b.낼�w�R�ma��[S�����P�B��!��B$"T�#Jr���� ��@�n}�
�ͻ�[
���H7AL�6o&�a��	� 4
_�u���}U�X�1ZM_)���h��P�|��z�= 7X���)�(B��471��2��
��@���'	�|�_?,�n�$����G�Q�Ir�����b~q��:R�οn|��B}���p�D}���,l��iU������7�>�+�),���� �����ߟ�\�E����\�8�����KN�L'���
����|/W����k1�C�6/� �O����^�/����e�V�q0%!a�Q?ּ��:�N��&{۰�j��>�vZ�]>�٬�Y1��Q��mr�`��������F�Pv#]�6� 5�Cv�"�����_��At���/d�SvY|L��O�{V�pR�W�}�^�ݥ{+���nyJ�F;�#�*�I�~��=��w%��L�ޒ�$1t����輢D�C�m�
��޵�u�ܿ̨�v4�L������+��FC1y6�����{&��ܟ[1b��Ս�^���~=a��*3��q��;c�g��ύ=�;�Cװ.�;��܍�D����"گz/���)n��G��ZP�[�/Z��`FI>7���K������}���`>���r��0�g �
2v��`.���B]�L�_gR:s�P��B�)���t��V�#�*X%��r`*sr��d���;�X�l,>%b�F�_�ś"3��&����h�g71��d,t{�����p+��x���,����+5�Mt�xWu�w�0�����H��)Me%5�Ȼ���D��F�1�b�s�T(�����h0�
:��4�M@��i���7d,��b5�u!����rג��}��'l��J�;-��i�|���3���B/T�}�J�n���˥.m�jn/�y��M��󥏿U4��v�ܤ�]0����q0��1��o>�w X�^b�����
�{-Q�`i.����H����Z�Z�0{�`�{{�Y�D��VҴo��W���a�s�Z=���������z�|�Őw�.��8�iA=�]�A9]����:��I�b�P���bA��/�$����4���l��yʳ-�2�̑Vٵ٠!���,��h[���V�kGtz�D�HL�؏L?�����|�񡴛-��@��JҳJ��mB�JƄ���c!n�[w��+i[qz�������1��	�nmdv֠w��|8qԨl�H_Ev�H`⣕ʭ��B1��R���Svm<*j	XE���&	� u�c�9r�Ûuג���eG��"��	��;i,^^�!PU$Ք�zNפ�K�����ɾ��eF�S��7�-���d�l<��J�[���c���s]ZKb�3��SL)q������t��B8^8R����Q�Sa�Ytf'���`��bqf�ɑ�/���(XH[�Uh����pZf��+-�l�
�g�;^���)�<��7$`1+T{9+��t�U�L����>r�́K%.	 P��9�K|�H��_&U 7�یԬNC��&�>� �<:����O�?,W��	�Ǥ*M�RvJ�̷\��{�Ų�i`�B��NU(Jz��/�qj�" ��ES5��pݺ9�����&�Q����C�8�e�op
�F��L5�wj8tq�mÏ@JTD|M ����������NHY%/�ԭ�l9ei�>#��W጗��X�mϲ.mZi��p��/��Y�lJ��5�i+���TP=֩ˬ�P��M
�xI!o�$uɧ��P��m���ٌzI��Qy��ŝB|PO6�	��!��C~�&��p������ۯR�"�_��s:�<�Ce�z��f�&��1��b�X!(Q04��\Z�#k� ��;D�_�F��~�.��/:��3M���:͹�\��PR�37ˈ�1����C���]��>�7�!���U&��Ϩ깐��hI�NG�$���0�D%-�5<�!0�_�RB�U
Y6z��O=��y=��N-�?�a�%O�בt[�-3�0w�\�d�I� ��P9�٤_�`�\Uea+�ӗ�!S�Ow1_/8��	�#���a�����ӣ�Z"cI�"��ג�#^�
�"}��Ju��T�����^��M���2�j}��#�c��B���������M���f�F�g�{\`r�è�ٳ�K�pr� � �/晴�U�jCh�aR�����e`D嫫����~WIK��w����@���Fb[k������)DsYB�j�U���$��1��/�ϸ�ֺ`P�zU��klc]L�J�J"���G_�EU�̔��q���Rk�,07���O�Y�[� k�D���B�0-C������bԃ�[+o{d���~.��i�۱�|�`���嗥S�� �T�@
�e�/R��S��{l�h���y2#�E�fƬ
��,����E�ۡ�ɥ'/I�2�a�~/��2'X�~���m��3q�e�w$�b��O,q�ŷ�}�U�{Z��2��U�����H%t�K_'���1��w2?�q,�����&e�B��Ƙ���H}|����ָ��t����>4��CTT��'�1��~���� ��bՠB>[p"e!R4�����������̣'��-��ߏ[;�'f���F˔�hɢ�����[��(Fb�JI1�����[�L�4L�D%��"�l@�&�!�'��a;�ue%��XY �ٚ�l�8��P�N����'�z)u�΂g���]�4^Av���4p6�����]+�*�k�)̘j
�G��O�y�^�<^�����Q��S|��|��O�b �կP��'���G��;&��a �D����S+~I�D�0h�M��F��y��Wd�8�s�08�xl�QI��&�2XF���T61�}�4^���q'�5��ӭ�$1��Z��@H���w��ېw�$������f��Xǒ���X�$F���O��T-�7_�Pb?���Ŗ����a�N^\x6\:�jT`A!����m�
�xL�c�ʵ�.v�vY��4��ms��a��v�e�χ׀� ��&%���cZ�����{h&�pB[�~x_W��a�W��o���|4��еC���j��t)awg��}{��k���4:L��z��tō;/�;�آ��g(�4��]<<M>��,D��~�$份,{��rp������r14��G��|��/����Z��Z&^o���#��\m8�C����h {�Ϲ ����LPT%�V���:���^�ĭ�
c��{�x.X��y=X�&�J �{I��Ϣ%aF��o�Lno:��g�#ﲳR�Jl?QqB�R�	���\HbuԪ2|'l7w�F�2ġ�B^Gi%n
Ý�f�_�V�"# �� �>��������\��?�v�����_�+�5���3���S��](T���P|�Ŋ^d�uxo!w����4�)Z�>�+�a�%�H=�
-��'4��

m�&گ�)���py�X�ihv+2����:�K֠��\2W��2�[w�� =Z���rDf~P��A^�9��¤�]���h?���XP9?= �F�T�킯�;u������� h���?g��"�0ʠ�)?tAn��
#�A7��v��m0��<�췥3�h�.�n�9��UF��J��
�".z������*�mmw�rL�D{*GC�:R��
�f��</J�8O�" �1R������rq��<D���Q8�������FW�~�P��no4�kq��M�۸!%��8�[��8�|T>�k�v_�� �@%��[����24	�U< �Y�"���5%+K:E�v����x��8)�nxE	���o�Iڑ��2I���j~�'�z��'�8�FpE��lx�Nǽ��I�{����=H^k��]�P+�b~�_�Ï8\��i	gߝ��>�k���V�ŗ@逴�W$��F��<�3äJ�WAU�k�5�;�'��h䲏*��Rj�����_T��,H���`�(�[�2Rٲ ���NO�W�[�6��,җ{�2/��7i�4��J(fԁ�dY w�{[�K2)?1p��;�d]�]I.as�����A��űtn�̉t��n���u�!��-�#fZ�6��s|��`֋���=GmyT�%	Im�􀐐$�F�f�\��� [*��������L��:��qL0�$%���4�`q"��#AA�!�{�|՞��)>�qǘ��N/hDg �H_����<
*�c)~d��j�p��PyB;MG(�jl�~���h�no}�,����ť�-��/|g6b��'z���c��R%���X��!m�8�67��xѕ�KJ�S�)����B+T�r`k�c6���e�/<�7��|9!xI�`ʗ�L�d�0H+q12sL�_�P,����Bꉅ�V\�E��x>9�|{$|�a��NҊ�~v�������&~�d} �*h�x��[�ɤ0u?j��LS�82�1�!\z�T�1?���5�"t�a �&rO4��~�7�~�`�ݘ������&1H"T4iEc��Q�]B��I��`�lL�����"�7�M���]q��\�s/���i+��*Tf�4�F�J�mk]9t9�IG�ސ��>�����{���s�rq�K DDu>�-Ɇ�d�ʸ�D�ô.��Ky�����b�s���i�3?��/BG�D�;����
��=�L�Ti�����S�U��e*Ç������[J�,�J�M��iָ�v�P��Zhu��.IE��M�\=�jm��������	�\��, H�vQ�_�.?[��	^�
�V��d���?��΃���PJ����k��V�<Y�(�3B.Ӯ���mv���߷�W<��ND�.���1�C���
��9����A.���&�W��Z�ɶBm�3���%��� Gl?���e�S9�����������nX�G`� ��(�R��P���M7BQZ{�@�L#�AE%�� :ׂ�����j�ivЩ�ٮL�D�9F�L�h�%[ٗ��^�c��l���!��o����r?#D	���Gh�k��'���ܝ��X���$�P�T$��Z)�i����~ڙ6F6�f��p�Mr�%�YX � Y���[9	��-۳W��Mg�NQ�@f�2��o���0T0^��p�$k���pI
r�D.����;�"���p:��-��ot��j�f%��b�m�n�k������~�J�b�-���5u,�Y�<�i^z��<t�%`ԫ��
���lg&L��+��C�d��Z��r��?��$Y̲]3��I�&�{���|dm k�I!R�fG�?�鴞0u����`z���'�k���� <��r��_��Q�"}�y-���N��[�]��&1���W�E���j�v���*��W���3�I�8{��R����: jX [�p�[S	˦�69p-YK���?��f���o���H(����!�	O"J��l�{j֮�gp�AO��Ӄ1�\!�X��С�d��V^�q
08p"�m���dѢ;�1A��i4$n�l�ȿ+�Cǻ�L�;'T�bA��P�M����~(_��[���aЬ�9�����Aڨ�j�jd>E�Ԓ���.r�	E@�;9����0	Z�窝31ʜs0�)���C���|ܪ�I;_��Cߖ쁌7e�B>���zjZ#�/��@�N�.k�#�v�AjτRm���Qid�Ȁ*t-�G�W����I�5��]̔