��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� rā�SZ )����C.��&0C]�-��[�3�-���+��պݣ�k�J�vo`�A�����f����u�X���v�=�а���]Q�Wۿ�߸�=_Q�X����j>��Zw�K��SvX��ƥ.���#�����Z�0���#7{��\S$��@1I�QX~TQ�E��db����۰� ���>0�%�9�j汈��}��1� ��2���h�G��SeY�a���	'<x�p��k�H`�H�j^y�0�s�78+���ֳ�`�R3dW��_��{p[�?$�s0��#�zS�_��bH
�c�p�IL7]� |����Q�� ��Rr���=��E즕2%�����`�^��l�q-�]�p��jf��Ӽ-f%H���ȳ�>��+���M�71��4_�) 3�46h�rb�J�W� k�h~K0�>P$�_n)���5�r�j��W�J&޴o��$>��6��ŀ�;A~<6P��K�~��f��*I
�Z��}`q���ApC��n���g���3��-�іrO�mF���,�$��@�BI�q�}��Ȥ֐����î�䂧��@������U���vU������ �T#K@f�㯁����|95<@���+�-�)�����K���FI�k���*@�m&���
���ma1[�2�u�I�\�U�yu���o�|��2����;�W�W�}P�K>%5�'�8���׫=����k��,�t�M�0�8]q3���N���GvZ�i�+ C�e
��Ќ�S�v<%���q��e_��
�k�夞��>ZO7E~��5k�TW Aod��eE���G���ɑ-'���?�G$����ќ����8ɸ+ 5ʗ���l�d��,�J�
�^�3b,�����J����#n�zK����z�&��;|�\�^���'e�W�����">�w*	FO�Δ��v���I�h�q׈�e0u[��E3�Ha���$���j�P��M����hvdR�\��F
[Y�h���f�w�jZ��Smy(��0w!�6�L����m��I��Ý��t-C���$�3��~L����o�Y�~΅:�`޺n�_Wn���'��Z���ZZu�q�;�k�3�J�[��m_��~���k݀�>>�Y�6�:�g"��9ZZP]�ť���st�6L�d2a@�0W������f�!(��ƮO>2�.�-.���̫MTw�RDg^O��},�oe!�����b,jLbX��|-��1�N��+a���h����ɊW���u�mC���A^��LPM�{���6�S��'�i��4���_,�B�d��AI<;0*��� D�O��˘@�����pB��h��-.f���	s�JpA"C��t~Bc4>�J�a5a����u[�V$�����A
��X3q� fv0|{}���=^��j���2{ r��G����1��;�:Q�$�qT-Vl�"i�y�}Z;��_0���,�hFhx��E���lS����ˇ�Q�O��F��|1�:Z��*�	=�/:b?G��gL������h�\g�I�h�u�(���&��h���4=rO���5�u�i�����-C}�\MJ�c~q�qbÏ׉Z:�g�H���lL1.GoϷ�g��Yi1kL�|�P��N��]>���+�f��9@"9���$��goN<:Y/��Q�(���w_M�����:���A��o�G������O���@��+`� z�3�����\��m��K�~g����An��v��Zݨ>U+���nS'n�Sz>�C?�������vIfI�[���w�j̦���W.����l��51gN�ZI#��K�v���<YjLD>(��[9쵿2r��Ņ����;Rt\�,{�o��;�d���g��
��[ZM���!�ϿU����XE�8�b�(��Fׯ��P<����eŜL�kل��nJ/5L�?3��G�-F����rp��NeVS\�����% �DDiV^��c��?o�T܀dh�J�ī�@ �
ܬGL2�h5)�	y�%�V��^��6�[M����&�\�(�nh8����T�}@�[�i&�tK�h�̈����_��,֕%'�/;�E���3pa�D��K�,-io:F��!_�t�-ƀ�3��s�`٢�-��	�$�oBRrY�i��K~��F=N��X��h�Z����Lb�R8=���}Eo�L��N�*���F�zq�a#��Ę3�юb3Ĵwu�z,m����i� �2�9��z^F��\oG��j�w��=��A�ӮG�����L[����.m]M�K�Y(s2�|d�jػ�4RI��M�R�*���:�3�a�}����&�����"L��fIS(��.M��E�>���Lv`ǥ���#g�k˽r6���be�&��r�p� _}_�����A�����3�h�/��~�ֳ�˅ZV�[�Yo���v�8VQΠ,�˽)�i�i��S��jND\��{!�]F@Y�B��Wc��j��+aE������w�.{��п��������J�z��]��2׈�y�du�C:8�렀U�If�Va�ݿ�w�?r�/���mღCs���.�d��و��̅�����I �V�tF��ε������0��8Ԯ��_>�:e"��p����7	�:����as���┙�vV0hV��e�MPa�z��E�┠U�a*����~�yG���F� ��c�c��7��V��Հ��!f��g�k	�+	уT3�ȗ�CP[�M���ަ�뷲�f
���E�؈�aљ���<��`r٠��Z(TvZ�dT��Rq8�a����ܖ��j�u�1����/&�DG8��#��Q��}��ԡ%�r��X�+��ƉS���S�(���?X5���6�ވ�g'�YHO���z�˕ڥrˣ�ܼ�k3F0(�j��~[��k��rL�R ����B��=
���F�N+��(�樒��r���.X�֮Y�u��6��2H�R��b.d8��	�_������AL�!Z�� �ߴ�6qw��p��Z�%�k@�i���sJ�z'����K��Ԙ^�������r��,d�G�ԉgy����Ǽ3��\P�ob�YiY �l���`����4:Z�HK�b�v�|Zn�yRn�[q�˕�����P�g��dԬq�H>I�L�� �	osf��*�3^��vt�s��V�*8��'�>�M]��PFC�'76��ɾ��8d2�Ľ�I��eA?�|�����y���MYj��cZYʐp"��3�lr�o�)	�а����MR2�L�����jɪ$?��8éUT�aI�~���
�F����wt:�5�;��>�=&�J��%���������v@�H'�VՎ_Dt37�F�-��k:N��)}'S�c�_NL���q��z�fDZEށ�:�3� h�7���Z����X;CsZᗮ@WM��i��m�=����5�$��D�Q�ܙ�n������
q�>>�ָ&6��A�ʽ#\�w������?�9x���SAc2����-�2�E;�"	�I �)�;rl��i2�`KmAcN��%8�Q�uRr�ґ����-	z#9ot"�.xsT'o�CC����|�T�d��b6��R6o�|y<Î�3�m���1��9
�|���bf��T��m���%�P:c�Ԧ!��T_=oȖ}�t�y�_��䮶�=����^e��f2���D�s	��p���A��]��o�����޼�usj�Pu'��g��|'v=8P6�+Ks1�����+���H��s�,iU�Sٌ���L�����,�0zG9l��� ;�C��N�S9�i��� E^ɰ�~�;\N�g�2��̢�Ѕ��c���vU�P?(g�<?��>0����e��H_�����|g���:�W1��J�ײ�R�����/i�F!��'��_n�*�\����D�F�䡉��3�$S6`�C��;H݅��bWZ�lN�~��!���;�|xx����Ը�ߚ�X̽.������.D-�{_T�����{xSR������ec_Q�j$�`�f*n.ɦ|�Q���+���e7e�?�S�uӽ��{%���f�FG~ּ��Ӟ���7i�g��d|���!~�=�S#R�Y>�uc�v�uJ�X:i!�l�QNm�	t����8��G�n5��?�6���/�'�*N����,�'�wl�ظ�HS�(��2�>d=���.:x{�Y���rwj�wл�H���m�ßO��B��&ZO&X3�p� �˩rT�S���1��q�]��tx�&*�����-��rP�|�&�8 F|*�N�^��_Y��/ꚠJ~s���S��^VtHF���Fy��jeK�?T���'U�Yh�s?����b�I�m���������-�bw�YH��㐑_�`�ѫ�E�;*<�jjWd�_�.J8�6�����0�S�M���Cd]�S�`��l�6B�?���I�1�[�����>����J@�VZ�ѕ�RT�o r��ɳ���3j�̦�rs�����{��l��l{��>XB_���?��#��n�܊.m�/�q��8t����Y�V�!��������p��f�64�Y�I���z��$�;�
��q#����9��A�s�@T`�bV(��(] tjSb^�C�?g��`�ǌ�KZ�N<Y�
��Dɠu9Jh�,�zBd��H�9��KuM9��Rq��c���fP�"�m�?�:I�P�Y��/�ޛ$:!ʹ'M�-�߸K(�@����L�������MU4�>?
f�e��������Ma�a�eg���4�����sTm�t�p����8S^Ec�e���L�a
|/}�ڗUf�W��u`���f�Z����T�:�I
ߍ&��"7��2��R#�a� 9Q��蕞���:E^o���S�@ҷ9�H��Q��ձ3_�&!;Ս�r�����q��L2ĥ�be&����/<u��ʹR���\�$?jaci��:c(W���6������(|fn��b��)�ZD�	p�����0U@oG�4��'B�T��r�]
�F���l����ģ�8���ƕ ��DY��[��TLoR��r���Q!��MhT-f�g������=��NvuF��r��Ci�Y�C0��$�7�Tg���v�ޡ�A#	U�~,O5�� A�k%]��m�yQv�5P񌧕�ĒZ���X�;����RQ�m�l�X�Ķ1Eް��HS�K�� �^��V�"��R3G�:�z
�L�A�ObX����b9��� G�L��X�6�[�]�E/��Ϊ=&8}�4��|�l���ڭOk�ΈM\��S!��u��h���Ԏp�Y��,M7�����͗���IB��U��q��;]oQ�ъ��.ڐ��i �UO"�K�{�<[m)u��_ϰ�_~KI��u�?z!ٮ&�xl%G�7,dS�3±28R�9t�4�3k(a��qV�a�T~.�>��ȹzB�;WQ���~6}�H�;��/��=�����#��)�����)at>]��Б�[Ρ�c_P�g�;�(��8j�ɷ}��$�u�`��H�ŵ<��a�G�ԡw�!���xԅh,z� ���W��$8��)�*�c�����6)D*��w�Y���C�q�����>���R��m*�}� ��`�R�s:#���Ųӂ�+��&�9�N����2y���IP&ˢ\���g���C�����#�Ĥ���/f3���r@�U�� .%��T ����w����d�Ś�U�iR[ɘy58f˲�-�����wQ1����hr�$�ac��l�dK���sD���f(:� A@������'DK���y���luzO�_�Rյ���}F���fM%� ���}4�s������g��N��Hk�:,�8!�~�_ꇋ9B�ަ�9S@���p�U@��DU�T�n���?kC�/�>UBΧ�U�~�!����Ŵ��'�Q����vjH*'�� ]$K�0��j����yZ���>;_��D�'^ ��{�l��c�������?�W;��P��rX��(�.��"��daG�l�]��>�q��S�[�;9��!Ⱦ�;�1U<�`����QY�(�������.VmlǦj����5�ɫ��߸�,�1���n�la��`?*����!�M\Γs�m��ݍ�7�4"|�#z�v��5R3�z�^��g]޼�t������9�w�/�����Pdn�T��Θ,��Ɍٽ�D�.uM!	jpN��ui"N�P ���ĻK�|7��E���ޡ����]5������
0d�����QN�Cߗ�`ѭٍ)�{_���$!����E4|�����J����uc�:������|C�&Ӱ�
f��.޿���Q�Y���'&�'��1~���b�M�@��%Mx;��$b]?���N�d�����x
�?J�Z��5��P&��uwv�LKk����5�JS���c��!<=��ͮ���~���QfjrK^
�ܟ�.&:�᤬�#�O�\g�r��T��ڗ2܆�G9Ʋ�ݖ�ah>k���@���"�Vr��I�Ο�� �G�p�[;l���$�ҭ�3��'î��V���i�}�x�C�w��$�������1�ս
S�yL�� 3���$���k]��0�C$ ۤ졙2C�_*�#���K�͑*���X�2�t���"�t&ƍ�H�E0`���xVa{}���`���0ӇS+�1��]�^� ���\^���U�:����>GMJ��4)�8i���9��������q��\ӺU*Ŝr��ĉҔ�2�h�Ԝ&��>|��j$��m{�u:���?����%�J�샟���V���U��BDT�L S!j�ɂ��[cx���9��_���4�=I*8�skU�.��d�Fg�'�"	{�U�N�B��ýA��H��0�j_�_P��u/���D�7���jK���h�K".ڼU���u�jQ��eO&�]��Z&/��. 2�%���r1<q��	����ca�`ab�ҟ�!��HU�,|��1�d�t-;��v�o֗9��Bg����%n�}��V����?f�sT+�6�u>����F���z��x�{NK�"C\o�i'�;�U?w���}Q���'�n�Y�Ǥ�e����}��K��[��.����/�u7S^fB�ݏe��.��jT��ˏC$2�沊���N�=¯�� ��9sdM�Ҵ�M�en��9�=(t�٤,�b��N���E���'�kw����h��������"S�D��j��-�}քlہ��3��s�|U�Z�OLRZ�<|�"�z�,�a2�:=���L�WK2�\�<ࣔ�e�m�.)~b*9L�?�c
�_�:&��tp4^F������̥�;���-�?\Qr!�J�c�[�+{9v�q$.XM�����17�:~��X����uebK?��mL�Q�P(�:��'n��U|��7�E!c��7y6�
�s��ӓ?��Ύ��5�M���fdPC�d�Ľ��EٱX���̢!�X@�@���������+��Axp����-���h�
2�
Uu��S����]7})�Q�K���+j's82��*�~\���׼f9QOVCea��6|$��W��mY/Z_UR膎y���p̗t5�`V��Ro,N�1�쭿��U�#i�0������Q�y�#��N�G��Ճ<̅��r�O�Նs�&3�})����{�7�S������U�gRb ޗ��A���'~45nUb�T]|�ꥍ�������x����3����;;�Ԝ��D7�x.V*�OLp���)Is�~�ң~�k`�{zB?�p!^�9���� i1��x� ���2��E@\�� ���/��1?I�ȬL8���/ǁ���������q[9�$1��]�
�Dӽ������ꪂ��ޑ��_?��g�%�L`$4����U�3H���ѐ��M�)���J�$Ly�ܞ�d����I��D�C�*q=���Ҷ SӼ>˵ģ�ZN�uG�����M����;��*F�؍l���[Z��������2��E��$`+�6�j �vI7v�5lY�ONr���t;�y|׆�ǒkB�۲���]�Xa��W�0
������V�<:U[5kle
�������~�I�_I`Q�����|-�l�#Q��}�����v6k�VAF}�Lj��͋�WKO���&��� �x�5E���	��ll\b ��'�m�>���\�ǣ/��[+�d9K�ʹq�K�n�"�1�����GP���`f�+�a-��COX��p@�z[��oP���q�Ix�ʩ��`0�X��#Z�`'$� �]�ݱ�vM��*4W��s:��q�+v�|�
{j��m@4���\���N�����ɶ8��p�s�¨M@���XdP����$�g}W��{+�ڒ6�^K8dxu�|x�����PV��9�k�2I�'ʉΠ�����I�V��;�8��W	Agˬvc���LF���&�O�]|�Iv�>GA0�Ԙ�.r�-��O!���3B��4025���`ӝ�+�k�Ɓ��G֩�Eo���� m����U�Yb47�n�>4��^ѿ������[p�?�]d�I�q�\N��@i�#��iT	L�č��`	= ��'�i���.=a���15�d����흔�O��9@ N�L��t�d�P��x�Kz@�ק����GN�@O���f*{.��2-�t.�>��:/^�jc�2LO��{��� ��4�b���b'X3�u1=�}b?���999�7�W!�9@���]$�u�2Z�����aEq=u���T������B����{���P�$�l�l��|X�|@?�B�v~E��+�1�M��l�k"Z�=��B2�R������1�.0)�_h�fVY����0�Y�?�-����8�چ��$�橉*T�١]�{�2����O��7��JY��^ �#�t�2�!O�m=qh����p�yR&��П�@d���1>å
�Yn��I>X� DrR ^f�1��8�+3�ow�Ӭ���I�Z�=NEH�g�3��yqs�%o�k�~��*/)��,���;j����ρ��?:�bkj�R�����8��	9P�ٷ�%���k�|��}�vZ��[5ۈ��X���LNc�R�ӑC�n�6�H/;6��b��׿�	�>�
������5�-Cz��%��v��i���{I���:@�%��_ݝ������I�}�u{��)�*�������aˆM�jC���=����d\+#�C9[�J?W'�D,/�W++3&R���߽f�\iY�����E�P����Fu
����S�``q֬tS��wd7���&���3Z����պD���$'\�¡\~z�s4?��I��M���"J$ Vd��a�3u0H�l̞i|Dl��v�՛>0�`ԝۖ�e��\I��	��N{�#�9�Q�=��	���4��{������[����;�����Wh�̳��Oo���}���v76�������)d��l/n��8x�VgN�;qF�M%Ē�>;���Ood��{���	}���1������M�٧�n�p��U�����r�z��xq I�^�R%g���Zb,�8_�6(r ���b(R3��/vq���.�����e����p�n�X�)��X_G�ӕR�`�xI��%ig�?�L=X�99�B�Kj�}���:�dg3��&�B}Ya��Uj���_䓩W�7.��}���BpiH<X��w�=99pL#�p�n������l��R#S�U��mC����1�Oa�h�9KgP��0*��b`Yr|T�m�u�C<��ZlOr8�yfPp`���qx�����DS�<��	vʑO���YN3G�#Ir''�&���3X�� ���ߖ�[��S�H�E3l�����g�2�*BJ�$;�����hC���/�5�m%�S����m\Ӹ��g5�m��_��`�+gzfl�cK\T,�q��8���s��yJ6�:��v�Ѭa��{Hʆ1���IƗ�X�&�!amd3�F ��"��dS���f�D�!�(�z��ȓ;ZO�@8 ��wx6�GN�EA?�'�\�jp��:x����\���8|�vI�V�(���^=���WD�c%Z��V�Bp9���B���~k@���(-��a)���h��۽^�G��Kn��S$��mVh�������1��x�ql Ug�;v{w�o�xh�څAT���ߓ���4l��B�,�1�Ԃ`������y��ZF8�9k�-Ǝ�Ϥ��=LPx._"�@j_��~F�pG˔�r+kM՗mp���
Kn�4ywt��lډ>�� o=�]rJ�B*T�_p�X�zi'>�\���PD=F��̥{�O�ʣ���|���]f�8sn6I����M�Cߝ	ɴ��
�+���5,���\o��k���P��cpZb��/�{�����"�gQ�$���+�_o���m�_:����6�Og�j�n��a�!�_��t�χn�ح�oq<aV=�fC�g�I��aĖ���˴R���|6��oZ�1;�=3X������!��z@�aw�|Jh��BV;��n� �O��̴ʙ�߆�:4[��=� }���<xޢ9���c���W�_�r��J<%{�Q�Ʊ|���eq�	�z�N;�V6��p*g�O~��?V^td��}w�����;(>������'BKE�vM�w�`6���	�M�I�Ao���������,���5�p�������a�_�܁�� �YpO�Ǻ.������%�8�|���@�l�d^��`�C�\��]�F�I����^Ӊ��)�>�a>$$���A3��C2�W���u�^Ob�էC5����$\Q�͐ME]�Q"I* \�W�j1NS��$�����.k`S�ƣf`8���I�?_4�C|2���[3u��y�L�R�3�^oxEVR�Vm���M�wIb�衖��p$�&�����'��bo�����y��">��Y����'Em��3��/p&=LC���d)��L�$�t%���B��Ȅ��^������W���~LJ�دp��oA!�ڮaHl~�C�*te5��l)*�g�6��J!,�|�T����}��D�U��AU�tj5��uͬ�6:����G+2���ľ��5E�9��&|!�,U���ň^�	z��$�AD^0c��>��ɳ�YN���.�V���������ő�pW��R섢���4E���Q��={
o:�k~�"����c�����:�Vٶ_�?��?�r�U��