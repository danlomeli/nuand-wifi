��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$��7�4��L+Q���+2�"H�������v�ao4��	�u��=��d=�>�iV�f��l0�Zs��7���~rM��U�`���e����K%�u��ݒ-� rā�SZ )����C.��&0C]�-��[�3�-���+��պݣ�k�J�vo`�A�����f����u�X���v�=�а���]Q�Wۿ�߸�=_Q�X����j>��Zw�K��SvX��ƥ.���#�����Z�0���#7{��\S$��@1I�QX~TQ�E��db����۰� ���>0�%�9�j汈��}��1� ��2���h�G��SeY�a���	'<x�p��k�H`�H�j^y�0�s�78+���ֳ�`�R3dW��_��{p[�?$�s0��#�zS�_��bH
�c�p�IL7]� |����Q�� ��Rr���=��E즕2%�����`�^��l�q-�]�p��jf��Ӽ-f%H���ȳ�>��+���M�71��4_�) 3�46h�rb�J�W� k�h~K0�>P$�_n)���5�r�j��W�J&޴o��$>��6��ŀ�;A~<6P��K�~��f��*I
�Z��}`q���ApC��n���g���3��-�іrO�mF���,�$��@�BI�q�}��Ȥ֐����î�䂧��@������U���vU������ �T#K@f�㯁����|95<@���+�-�)�����K���FI�k���*@�m&���
���ma1[�2�u�I�\�U�yu���o�|��2����;�W�W�}P�K>%5�'�8���׫=����k��,�t�M�0�8]q3���N���GvZ�i�+ C�e
��Ќ�S�v<%���q��e_��
�k�夞��>ZO7E~��5k�TW Aod��eE���G���ɑ��f��	��&�o6�[������9��]�E>��iR�P<�htۘ�B��ʟJ2{/;���`x!�hX!��ii�='�РO.���g�~/�ި��!�/K
!�9��X�V����H�`<�{��
j�Z|�Q�RA�H��<�J������C��N �`��W�Hb��9�\�H".'���2�:)B�վ�8���Xﮗ�3��+>�G�	��Z#����~;$t��{;��T.[��R>/����e��*�&H�-�tġOR~q���x�����*"��<U�p��h�L�E���@�t�ے�w��0���)+�u��q�O��q��݉G���� 0U���pgR�����sQ}�D�����
:0����]��\��n_�q�1���'�HB٩Z)U�&�6�����b�>V� &��t�Ӂ*]���&@��9֗��?�����%�{��;���PN'��!Jǝ�A��1�P�gO�cE�\���B,�wu�e�-M �=D��\�#��=g ��z�/#u)i��s�����;�xI|hA$pt��ɑ�	��Jm8�:�.6��z�C~���r�����4Zȑ��L�r�Y	K妘F(I�}�	h�ъ�:�ο�mI�|��/)��Dr�w�2(w����HB�k�Y���{2Z��X�3��4Ѷ�2���U�!��a×y�����N�/ǉ.7GT[3�u}?�w���	�U�)� ����'�1 Z�D����_�q�(��+�r�n@������+� �Pے�κ� ڙ��>��P��Z�)�0_���D&������W-�6���ja7���}�S"�Y$�wUB����l~�3���U<;��B��@:�gKK�E�r��=�����G�M��P�Bp����I�웬�)�3���B��v�R���p�6;^�6,ꀣuP{
��I�߶ǹ�):��)��by�"�DrJO�U&`��N;�z��:�a����k�����+p���Z�>��D����<r����l;�+}F�u� �tgW�j�U��=wҽ��ړ�8�e�����ūoLB�Yxx�⭉��@�[8��۶��lnH���l��j�h��JUF��MJ�z�y�v��rRnB���7�VDi��+\�}��P6�풃?Gh�x��Ew.j�ڟ������;.�v�U��}���À�6���,g�J�@r�旬k���s-^n:q�D��r2��Z���8pp��M%��^uq=���=HB֓���۟c_m��<�����|>��g;8:��=8�l�������'�E���sȊ������"��¶~
��C[X�9�<��;@�TJzïYB{8A���ӎwi7H��M�:PO�����������$}Zr��&�W�G�����g^���7���I�0��"�NP�+�I$)>k4�{�.y��} ��8�F�'��/H_kZ���fD.~�!L�aFj�U�@1�uD����W�'N���"���P۪L
�E^zH�:B.�c�c�K;��l��.�$��S��p ��v�/���^�nL�K��:K�B����O�l�⮔a���LP%*^����ّ�4����z�WW� 9A�چF�̂�v{X���5��[��C3 4s�����v���)�O��\6l^�=���^O�H�p�d8^�z0f������*�߆g�}˲y������!�L߬��xV���S�[��b�X�Kl�o��;�pSo��_W�Dt��y����D�l��|�FJ�t�܏�sc3�^��;SA}��T�\"j�r�������Jlz���#�� :C�'b�!�$b�_�J���괫&Ԯ���y&NUPߋ�����g��š�v�� 	7��vx�"E�������OT��?�V����q��чEG�r��}5#v1�m�����Ex�^�Ǒ�c�=r�`\��9#13�k�I��sR�w4����@'�K-s��
�j���E���DS������(ۑ�tR��5BI:��<��^˦�i�!.Z�� Q)���uo�p�&��"o?-�(�Ԝ��B��gb1%`�aKY�XB�I�	�a��5�`��|`��G?�e�F��t[���qq�o�2������Ex��a�H��W
ZHq��G!�ċi���H�c�NױWȁ�K��a�~���Ѱ�i��[���{�G�Q�r��쳞R1�<}F�/ʗ����}G�D�F�p/��"�w\4noK�ߙ����\+"�\"N
�
�&b��~5��l F���V%��NkY���ɀq�z���sm�$Ⱥ�8�K�u���~���d#G�O�ȣ����}j�j�҇g�D|4�#�>P�S��W�	Ǝ6s�
F�gm�yh� ��� `�@#{�O�];Ia�r�� �Pдp���p�/��]%��.Z�϶ܔ#�L�c��?O�T<rF�S�]�@�?r���E������5v�:^U�H���M%����_C]���Ak�(�kk�'c��bД݄ܺ6]�L����K�EP��k$��6Yӎ��6kNF|z���:��)�x"4B�L (1�2Y\N�(g@ʽ�)���'���ev�T�Ou"��GGS>�~]�&m�%?(�f)2N0Ǣt�����dƚ�����J��jy�}#����m�[n����W���J��:��?*O
���=��x/,V��	c�����A��M��j\��I��F}mM����>���jȫo�~�qպ�6 6� �Y"z�h;N<5I��$e�!�4b}H/�7Ǉ򤚘�jE7𿙬n�};%���I�C�G�o�Nr����m�5?�"k����a$�7����o�~t�;E�P$����7(;�roa�k��?`��G���)�n2a���!*�2�N^f�'��ߛt{V�%��f-�v�ewvrdh��+(�����!���~��N�Ա�O��;��f^���5���+ym��H��}�1��I쇲lٶ���Nhw���qĲ\�q���ؒ��2��͋6+�|��w#LW�3��#T9��s��?��a�#�@��.7P�t���(���D�q���&�}�s�S#�:�-, ��~�_O�NO<LH@6�1^�j���	���T`�ֹs^�*��x�i��/z(�؏E��X|
Y�*�_M
s
bGB���IY���$�!3!ź�#�HzbRB��0WN�H5���W�R��|��Yܵ_�PR�B�?�Я��$=��2JqF��P�GJȤC�]����Y2���7���<�c=��|��8�g;�������7~��7�\�D&K�`C�B"�`C�,�����.���`K�S<x�/�w�̶pï����D�N�p�����O����!��A�9r�	����&�b�,�!�(�*��nFڣ1�LT�i��/PdcC"R�G�V�g��D�]���vRm�SW��`)X���B����&
������I�'���;����k���))?�Jc��*���ȫ+&T�A2���_*����ב��R���� |m��0:���P}�yZ�
�_X�b�"3g�+��;�VF�qV�����Ynl��]V�guM!b�,<��5����t-��n>\J��0v�,#��})�U}����>*0X�#��a�!�EU����t0�2��Q��,q�+v�/"�a����c��:�BY;����)�RK0��W���:�Y�}��|c�;�;�M|A�&|1�]�X'��y?\�J�B"�"���Y}�cRh<ǡ]S������?h�`��zJ^Ld��6���T��ܽط	Lت����y�m>;��f����$�>��m{  �����W�Jv�3*4L�ϸY\��F�����������l�G�Ͽ�Zٱs�� �(xq9.����(��k ��r���u�o3e*,Y`�zP= 3�ȡ+�~��Ii�'�dd�����*�b�9H�����9��!�]�Qm�Oy��&��	P�}NH�F]�J&�i��	R���l��	*��pp�*�#���a<��$�0O
.ݬ3՛$(ԃ�(����%�=�����5�I��Y�%PB�ʳ�[�C�,Jo,ї�Hp�9.=��=��L���L�%/8�H�{�f�\0������sت��I(VU�bjX��L�ђ���:�&i�y��Eޗ�
+E���r�w(����v,nB��>}��~ɞ# �I��u}�9q<���T��]P�|�m�@��6k��Xw)<�k��[KxH����7�NZ����L��١Uqfn���xW�Zb�e�p�x�,Ѭ��-�v� �Λ���I��	��T#�X��4��
�4��I�6)� 7{�VȀ	کY\�+:s}��ԗ���������J���wDO��ʩ���d�3"����6�y��{�SLM��c��}C�Ï%d;�q��
p��?�ط٧��G���+Ф�p6�\>��+|��1�r��<�a���.�l��O��4F����Ld��h��|�E�}V�`��YR.��(���·",	[�-3�]o���H��]>rT�R7��\i��*��e���i�m>��8I����5	��{LL�`˕��0\���6�n�ɍˉ���W�;ɊǞ�[#-�Iˡ���/����O��e���'��X�b��W����Q����iTlĭ.0�s���U$�bF��w=��r�$h�������!��I���z�?B�����D�f� ���L�}�¶��"X�WE�����q����ΰ"I� 4XPN��Ei���*F�w^x��������>y����O����ֽs����ˮj���[�݁U��ܪ���k�E��p��b%�ȇ�x��*w3�Z��N3nN�>�Kw�*b~~�ϴ#�����.K�9J���8����B�,�!����G9��w�JZ13��P����[s0B
��R���,�����5p�k������Z��KVB:���fM<���Y��d�@8ȇʍ��齁�c0�w����z%���W���z/�N��`L��R$٠ݬ���#�x��&H߫ԛ_�����J�*"-�qG���)ޝn��Q<�q"�w����t��KM��r���$M�z'�7�Bl�[�ډ�E2ly1��Vej��������OI�*�E���w6Q�C+>���[g8.����i7�L��aQ���m1�>����H]��F�(_A�_7a���Ό���B����g1���t��;T�{Qsi�Wo��m¥���:��DZ�.Eq�A���v��$.��_fG&3{+�veW��Y�M�l�9�h3��'�<9���=��t��{�Т�Mkm�iN8 ~EQ,f:1���F�.����>m�l��d�M�0�o~A�ak��VU�%��p��|�䒑eXV�)bJ��֨�*	���_y��n��6��� �J� ��l_;�{<�%��� B�����3(N��!�ye�ȿ���Y���k~s�	�� �<�O;���S�ܳ���'�Z�H�����Ė�Ip5�;J����m��±��A�f-9���	�k�.�Z-fʗ�˝r)v��Sovw���s$J#_�Jz�)�ԫ#z������O�'悮N+�c��Ͱ=�x��)���S��,`S�ņ��hU�s7��xGY��#�9+��>��� ���v�珝�K�G�j�x?KEE����S<�tK���ze? c���vvn������j@+�L�x]޶�6$8�9�;b�/����DY��G��01�Kڲb�k�;������2��U�78���[��L{ܹ�����8���HLf?,a��4�7q(��`g�M�R
������Ʒ��W�%��x����/ǭ�۔�:�@p&��l�eNЇ�ld h���=��&��S_2#:_@�w�u�Z��5IYkt��1�'ej?�>�/�=0}�aU�����5káCaQX��*��m����ؑ�,?�cc�	�@)[�����شr��n~]�ю��Q�C�� ,��`@.�ЬC�ߐ#�Ш�	����*ΕRռ���;)���=x�N˞M��3�g�~`�a��P�ٺq�D�-�c2�Ho�P��2����c-�,3�h��/"�?6E��D�+�/��0�����͙�j����*I�f����*�QETz�y��n��܇d9� a� �7;�2�I�Sʼ)ɤ�����n�	N�c��þ����M�du��͖�;=�������-Iwm�\le a�l�v`���g�]�v[D�K��P�B�{%0�˚�l���܄N>���P���8�Ic_�z	�p�^�
�i4��;�[�`�S'��e(Ğ��*��٤��q^�l<�e��Ut��$�hǓ���"��eS]��M��]8�#I�#���m��V���i�s����rX&����h�4�����%kg>�V�O��j�(�x�P���M��i�g�����n-�9�;$�ᓡn�0�͇�Ca���SS��-�T��]�d.�~\n�V d3��A��/!�|J�)�P1H�щ�"�f���J\��K8����V��xآ˂�V�.�A/X�yDL#� ��k�-�D��.S�`��9����`M�u�9�R��a��\`�7��[�U�&�P�(�>�{}��^���Z~�c}Q(X�	��o�hp��Vb��6^	�_�5Tz�S�	���cg+޻i��͹�	X;5���6����]�����/Љ��JyxI�����g.��?$��P��i��s�$H���@���S���c���a��)BT/(q)8w���T���zWi�����SB'.�'f2p9�k`�{��y�a�M$�8J�b�NSԫ��TPU��0)�����D~��Fu�; *�ޱ��S(ZF����ϕ�y[t��&pf�ibXx&��0o��\��z��A-�A��3�_����) ���sR���I���Ww�V��	���`ȕ�/ɵ�{���x�ܭ3�:3���#�X�+�hz^�����7�C�1��lZ	t}�5d�,�p��ϲ��%p�=�� �˄��_oYqr�[���X�֦X�L~.���)�Z8��+l��ȴ�����RӘ�P�K �zt�vAU�]�D�4"�:'qk,� ��T�L��e�.j�nXX���/�c�M���W�x���
���+.��M/�$��z���S��(%"Ԡ�9�8�DZ��fm�#J� ���x����a���~ ��Ԋ�c�=*��*ܥ�����xQ�N��s���*_�Vd���.�����FE6���I=��{��wi�B�y� �˸� ��v5q�]B.�Y�u~� �݂Q�6\'gzAl ���i�d<�z���~ճ���=��v'��C�a�@W���FZ���xCq7��!�AK��v�gF�Y$7�;ծ��7_��E��M���'WA�I|�	#F����=�;����_ �{��'=Mӭ�e||�&��#-N�2����D�6J9�YXjE�Ґ��[��XB_<A�[y�sMC[A�&$��1)��t�{J�8�ΨM��X%�����ŴOWy��Vcq��Ɛm�(.@��N��l�>�M0t��B��.[�m~�~��ػ }%���{�z��YJ��J!��j���KvJnI�B�@$`
>TXK3�j�������<"�(y�����į�\h"!���/�Vb*`�m�n݄�xF�h���"k�R&71,�[�p"��������W.�e��[��Įy��>ۉ�p�"]���˼l�y��M�#пe[���eZD�wWZ'��v�8H3~yݶ�U�bΈ!C}y�`�Zn {���e(}X
y�V������ȥ�m�v�y������vd"���J� �5�9Y��1?7 ��MN������2(c��n���n������_�%�E��\��_?�$$�a�����g{���u��7�D�Q��@� �?�m�\�A�@pC��b����Q|ܲ�α���R_`ږ�k����I�u��t���^�3��s����5,�}7��?e�&I{��r��!"�G�0����J}�G�/Uk�\h����qd�4�;�$�?��SK���M�7���R&H �6�R�i��ac�sg�H
�@��b�V|�2'̕)y����KӃ�q`N����9�� ��Fu���oĕq*yZ\�{� �R:�J �*� ��o��.�YDL��=݉������GY���ӻ�{�b�.�d��wn�L<Ɨi�4Xl�����I��_Hp)�"\�M�=��v����eD�O���u��]H�	��ԋ�Ԣ.��g
u���#Iefv�?�|K�+D\���!pz�梴�2�Yn�Ջ�Ȳ�{'h�~_�� vtB�B�E�Xp�|��@1�e]���GMZ �[y�E]@�P���E�l!��{
D���e[��԰�p��]"%CW��PN���rd=��D#"]V%��a�D��?�x+��u7�H>^�(���~�����l��iy�� 4R��W}��xfk�@H���uvT��up��)=�f��Q*��5���� �MƂ^���Rm��u�ɻ*1�h�"�ᘰ�?o�ˬ �}		��x���Z��͠ۍa�JK�n���(<c��*_�.�v��r�ϫuo-�	'��1�`���e����Nx82��x��]%3�%= ��A$iG�]�L�`���(lK��M��K�_�Dk?�.n7��Ǔ�w��� �*D9��ԭc�V���jۏB`�k�F�����i�9��ZΩ��2s�t�����pף!\��qd���VP�Qg�0ڧ��F���Q��{�f]W����W������Y��2��
D�_Z&/\^@I�O��U9�QP�����{�}�Xw�������d�w��]�%�����%V���(dg�M3�����g�%;�{����
 ^/���c�����T¤mvm=�N)Y���$L�o�p+4X��+�Gu=�g�.K�B������'��]4�5��sz�'W�-zu�I�6S)��W p��5��pF�����)c�`�󒟰�����G��)�\r$U�;�����|_)�)bd�%$#��r�6y�t&��ӓP�mZ���3-Ds[a��b���G�� �����x�����.^X��d{P�/w�uz/�Aag��+���sۛ�a,�S��Z�m��d�3���z�����KN�4��p�p�����Q�O�5����:��F���2�]���yNY.7��t���R���\������ � ,M�o��Oz	O��mδ���%>�� B����C���e��"�0Ƅ�`��S^3���3/���2�b��j�0��r,��(�d�`Pܳ�6MŮ������0��B$�Sҏ������:}p�Ga�=�6�� �He�]\Qr�pN,O��g�O�ܳ�wW����sd�[��4���.��cM���!et/XX15<�BR��.Hm���
�=�}�f��L�Fݹt��Z��v�"x2�m�T�\�	��W>BҤiN��Ύ��G�$9md���O�Z�1F �LՂ���)��Hԝ��:i�E�T+_� ��uqe��v/�ڽ���6���nN�~����F �����_�ҿbT��qN���O��ۡ;䤨:�#8����_�������yN�H0�F�3�����ҙ8���k�����/-�v���.Ha�z9����=��Ŕ�x�D.C���R:�v:��%z��`�Pq�bH�f�L��7v��&�(�����N�bBƘ>�Qx_%`82���¯��zЂ	��z��dҰ��5�p�
�Ol2yZ��b���@����% z��1Ԣ)����uPwQ�"NP�}.�i.��)��2�_D��1�Pn�(L����+/��BQ^�?��])rcQ}��~즕�\0���3ܪ�Ѩn�As\�vw������G�mm&w�,���G|D�e�������Ț�KO5� 
��}8���^\�����b;�W�gK=���b�U����\��a|?��9:M�ڶ-�S����I��u\���Ɛ���o�9WE`o���~IG����[C��AQ��c�s;���-NrS�#JJT"z�Լ*��c����/$��)H�X2���La��(!�l��P�ŧdV�� h"�U��$���d��E��zBE����_ QC��~\��%d�3ȏx4=J8+#q�����L�2�'l)���׆���'_��Y�0'/L�Og��+E����F=�e�	5h�u~�1|0ؠaB��	%h)[pn{E���My�ҿ��7�0�(�t��ѕ�^8��&;����T�<��;t�t~��Lk�P�RW~ǖ��8_{��]p*.�K2H坢x��,���f�Ѽ���۸I���4���\��Jf1�`"mʶ�,2����R��7���W�����DT���a�~[�w���N�0 ����ɣ핔�E!~�(�x�_ڰ2���3�
0�P�����(V�V�3��]����Ίa8
= ���T�;	�L���d�wK��U��B�3�p��Q�1%R[R æJ�Z� �F�j�vE'R Ϋ�F%��j�>�*��K�+��rF��ʁ��J>�3���A׶no�g�:"D��Ǉ'�`%q�|4Y��^��ȬW�H��[��[�`��
,}��}sA8#�5K+��&!L4懭-�<�/��&�um����d
q��w����(N�;��"0��E�wd�{���v��[5�5���a�ꞥ���I��G����ր�G�:�hufeia���#�8i4r.\"`��u�;�ݾ�߯�s���Bs�VΪKv�]ӌd���DfpF<z�����+���o�|O&�����.y��"%4&�n����=�����; T�0}X0��H��9�.�ѱݗ���������^&��n�eѨ����;�Ђ���1��+G|�5n�\�}�}Y%�}����X�U�7�p���{Rm�
-���{�x���T����R��%L@�K��R��^�'�fW�_��H[� v&����!i8Y�����.>�� �=��E����8J&�ԣ�\�4�#dCUv�M��J9|sr2���9V�;@+�]��7 �,1�r�~��A����q(��n��ڪߒ�y溊7��gE�9�h�i� �aJ��:r��]�P���]V��Q"]�^ޤ�-��,� G���w#98#�*�h%�5>��+	h��6����F����m��ď'�6��s���O-
m��[�A����s[#�#'�3�?�ܟKn:??�W�*��U(Սo)r07�3h>,{T4�ۂi:.����6������3yu����ݦݺ 9���H�Gc�� ��]�gU�f�s
�X���X��	�Ɇ	�* ��vȆ���V&��A�����t��/$F��S��8	����Z��_���.�6�:B�x'�=T��d�tp�a�C}��
�`4{�E���h厲*�iTh,sx�_��ϕ�Pׇ����&F!�����Mh�����Ґ�~�@���A��PĚ�;Z�� S����k�C�r�o�m�і�lj�o>i|-#����?��d�$5r$�W�*��GD�8�tS�(M�Z���+u\�<����9X��r��=��M|�۷�	��1âmtpj�G�e	c}
��>����G������\h�f3H��lf_O�wݸ�N{]�9H6��]7��c0`n?���C�����:��.朢��9�ꆹ^*��f�mdӏ���L3����9��<���H-��߹tct�B5�<�Y+,��TQ�`�4?��e�Q��A�:,��S��(�e����(�)w+���)zL��M��w�&��|C��Ǫ�^�X�O���+@�9N�Z� �rAr�F�+�k��Q0�3��X�.U
��N
��aHf��C;/�ދ�*=���!��6. �b��h��w���S�[ť����[|'ؤ����G8�� �%dʐS$�\�>�3��:����^�-�zIZ���,��4�$+~T3l�,L�Ծ�y����#+�mqc3T�����Ag;Q.D�.����Ά�s�������Z|��Ѹ�����F��� :ν.�l�I���S�Q�,?������m��6Nь�<ib��NW٣xj��9���ڗTG�qh����-�����u]������'��}ĦJй��4k������'�FE���`5��̈́2+徭}h#�t\�'n��Ѫ��W��_'�|/|�V�����J�h�AK����!nꔢf���p�1:��6��z1#O��#Õ�aYl�D|�}رY�Wss����=J�|�WƔ�����Ҭ���}���?���t�h��'�6-%� �U�p�?2ԩJL~Yᗭ�#�5ˤ�`�$�D��@gՠ4-A��|�y�G���u�*�������vyo[%,T�/��^�A�\�˽�-��h�m>�xC��!���!�����.�gӑL�w\�%�,c�L�5T������q�˘�C3���s�w@٬o�����A")�@�I��[y�h
�#쪽�8��E�������t$�$�T�{�g�MK:3���e�b1�F�� �Q�PuHu+�π`��rQ��=��.xV�3ԕgSc�v�����a���;��L$�6x��D��t��)���,ƉNV���U�1"��d�TL�NN�]m
�D�|#S�f��A��p�gZ啛i���_���5�?��b�k����P|�ӯ-��eKFɦ6xJzd�hk���.��[���H��c����!��ڻq�����{!������\�%�$:Y�����g�w�,MN���c�'#B�؜���`�ԷX�[�n%"���x͸����lߍ�VK�r�~.�4/�j��<S��_bz�X=���}i�]#|�xD����QC�܁ݱ��GDPm')r�p$�!�v��$)j�I��<�r/ʐ����̟`X��CqmҖ `�f��oް�>+�ۨ̽���ك>ɱa�hdi�X��.I�F�jR`�G����i�k�/O-�0�Z��*���=��(?kW%��3���6������xs;4��t�Le��)s��{�0�	��ΊG��ZU� zJ��8�S��z��j_��lN�Q�9��?I�w�U�N{9����*L�=��)$�ٹ��a0}�� �w�i�3\W��1Ww����}(�Ӂ�K�����	�����)���S��(���~	�W�U��p'�f�m��֐��#i�(�²^� ZC�`���.-�1zi]ȉE���+�xu�"^��Q��o�"��EUDH,Ղ�@ҷ���R��V�����`^���p�z9��p�,�����{��z�`ڞ�>䬰
�"��!�kd(4��X�f����T٫�[��(2�m�l6�̇�����[��]� ���@�8.��p�Ή=�xf晫Z�&�<����u�3Z���b 5C�p6��:ŕ���t�������U=iИ6a���lm<�_PgGT/~`|�e�^����.M�nߨ�P�Σ�Z�L�#�1�㓑�E�8�,l���WC~�!K���!O�Ho�*$z\���l!}����+��k�휷i7�:�3�o�Pq�_� �T����ԫ�D�+�>�[���������� g���*���Y�'��!�D��&]ҊSrP�>٢������c�������hL"��	x�'#aZ�'�z�,���H�Ia��v2!��]˚��V#�H��-�l�8\���sFB,闈�[���Z�A���LZT�uog�������aa�~O�̕!:y�>^��r�ܜ"RZy#��'<�tl��>�&�ð����$i�eo��Z��N��p�/Ė�m�	}�%w-�U"K��N�ε(���Q����ɠ��k���U���T���G�ބR�d&��/W�(CU��VT�Lka���h^e^��=)��I�|�[R�̽wN�I�Z��*�z��6�V�"�&�2/eN��(�7�C��X���?ĸ�]��/��Ha�C�!_H�����Ek�iL&@^{Mh})-��Y��5���n1��R���;��A��A-�*;�pqN3v�8gR�K.�X����5�G��=�Nk�P $G����+g&�(����{}d�!Ԃ�A�ǈ�ʗz����6&��KC*s��:�
͑׿�%��=Q1�W>+��u
`}�{�)]�HQdc&�=�A��[o�s�=?҈PG 7��g���k�Q�:�ϊ���Y:|���j��W(c��,�	.�Xt�f�����Uk�j��%���B�QӪ%1	""ܷ�qL��M����{�6�}l[Zk�֘�S���S�0,��)O�� �_��熕$86r.�d]\�?i�b�߅�Jk�<~���6b�bws��p��hԨ�`��+2�>��Yr:ĕ�$C4���i4���ؾ~���dX�ʨ���&Z�&1xReMl�[ ��vAT��$���b?�jW7L6�+���Ep|��>#Hl���rIu���q]5�w"h1�1�U�]!�Z	-�:2wAn?�^�2�3*!��y� �3�$P%X�8C翝&��]�&�l���P.�6��b6-v7�y��L*�"�v/�3:i۪`J�N�l
��|�͆��r1�0/�Q��TGv$�ÿ?�K�@�a�ʁ&��R�I2�{De,q������r��U��2�Y�h����l*�{���]WDu|J������|ْ�E�����!�%	L��09W�HB���*���Iς�V_R
�<��}��Vh��<��\B�xLЇ�(3����Cf���;s%0�
�N'��V���N@L��}c���5��G��.~�C�1�=��~�8�I�����b�k�fZ����F�� ��Ґgi�tW�N?{$L ��E�=B6����w\��>��dB�N.	J�x��S[�I>�܃=����,�A=2���:��M.5�/����Ӝ�
sAJ�i"3��Y���b].�>A��r���"��d|k���kE�tҎZ�K��˷^����#2\p
m��f��C��m���%@�������g*.s�c�r���	��Ň��.x�ʉ��93��I��|�;4?�)9[�n�h��y7-���Z"��U�r�p5�DF�#9@�΁��r��BnB�("�C�`���5*T?q74�D"��A9z�h��p����L������^Q�����\QQ�?�'��7�D�aZ4i�m���$[�+��qǨ�p=� �w��� ~1�I���?�ө�������&�J����T��p�N�Ȁ}E�RNm�w��r���o�LĘ0��"���y<�(����g^e|ϓ�$�Pv��@�SwMn���JY��#�kS�D٤Mv�[��p�-�>�^�	˦�!�����J)�`�!�/����U��KE�li��!�W����d:��ܝ:���M8����Xh�F�O3��Wf����}RA2��N�]���}ZЇ��N�> H���`�t?5=�.Ĺ�|�����n�y�&����U�7���ߍ��x����<'�pF�#Np���p���~����Wg��z գw��{̄�M[ujݳr����h.C�V")Yݺݪh�Y����M�!����%򆭲2H���X�[��u�e�7����$,{s�Cs�8��P�?��GF�:�1����͊6c�@�	$B�%�������<�Q�ȍ'B&3���ڕ���_<6�x�m��⊻w�DvsG]�]��|�%П>���[��c��L������3�"4�7v��2��|o�{s�In�����Gy7w�1���
�RJ��78����R�4�b�0z����e�c˶>(�1հ�D+�J���ʦfn�L�t�%`�;x�I��WT	��\6�\�ϳR��=6q(�O:��&�k�Ӽ|��ւTR��Ã����h�BH���r^�6�P�]�(�G�Vұ,�o���49�г�qôoS$S��0�3p�o΃����c�,���7n<��I����@`>�D���	�bOV�ҕ�l���"���Oo��g�o-V*��y�қ�"��egpV"�����2mUƯE�S�,�/:E��ce­]�X��]q�gD"�F緿���;��D�VoIݻ��.��bME5��X���)�r���),�5�1��-���)�7gb�Ѧ������d�J�c�����#.�|"%X��o�1:ymPgs*U�|X�Q��'r�+��^~)P5`x�,_rJ������	�ؼB�/��N^'\��	e�砪���x�>k����d�J��`,5<�&�p#�,�%�ĸ�g8}|����F��f	��;|=l�I4�k�x�9%��d��
�V]�7�$<�,}/���X�3���t�=��f�k<��u�v#��`f��9��M����}�t�ʾ4ۀ��(�(�;!�Ӱ��[4�#����sM��nۧ��L��j���Y-��e����AT&r3��	�W�(���ۯI} ��a��n��^(�2��l'/���C����4�OB)��
��0Ӑ5E�N�M�y��4:����(�?*8�$���4An���ʏ���7;Wh���h'�t
��[�*�ʇ}���wZ�It�e�KD��J_)td���/�.z*�&���S�o#0��߳Ų�6gƬg!/t���� ��.��ڳ��im�MHe���`���m��[���B6~��ʰUH����q�>��m���*1����	�`x����g��6�3��<���W�x�����Ϝ{���5�K���;E�^��H��E��u�i�ײ�2A�J��_69S��k'��=��ˆ�S|
��ȷi'�}��*d��MG<�����O	��Q���Q���G ]�v%��K���G�����,�M
��Ϡ���&p5�&�R����D�[�SW��Ó���Y�e
p��I >����3��j�ZP�HA�Ξ����3��d&�O���{E�U;�K��;�6�6r��n}J!^���fWH��AO��[�������Y��/6�h����T�Rmq_R`���Mc����H�ZTX�������؊��>(A8�w��xέ	(�����qW3��Ն���:�c���65��H,�ud>$��A3�XX^6l�i��� F��\R'����%
�bFg����T�b"`DW��F�e +�V�B�m.NF;�E����*Dyț�F�v��@Ə%9<������j+d��ۍ�
 ���@#�z��@,J��{T�v�~5ӌ��-�'�V$��Jr/����SO>�(�Ս��t��SPZ|p%��N2h�,:���KV��}s���"d�E_��pR�v��ފ���}���#��S�%!���W��7Z��ޯ����?�Q�Q�~S9_�ڍ.�,�+����Y�l��Z�/��>�W�]rI�ъ�3��^ˈg�=oM���q7ٰ�)v�q��V��Y�n�|~�.�����M�g"H�#�^<0����
#���w>��]�����7���pqK�lDO��:`��Uۣv�Zl���]:�x�њ��Rէ�
��-aƯNP���EZ�Rq�&�B�>��m�b�Q���w�P�t.�����y���>�s~sM��;��!^r����?_(i �T{���J��3;��t�)�+H���H�L~���1ɰ
�(2���m-9>��o�J����^�#��V	Q���A��6s��H����D웺FĬ>n�PG�f (vӐ?"/��{h�ң�(���sT3
X�X��azb�0З��çD�k ��icm2/h
�*�|�{�h�.U2q���Y*�^��Uˢ�ro�iHU�|VE�tԫ��<r[l�ϽHe����lӧэ��UuOE\dqaр����z���Z=���9��re�?�>a (:�
uV�Y��ѵ_|ӡZ3G|��G���*�R_:�����7���=~�5'n��.����k����iө�	I� E��]�%K�����[[�4-�#�M�DY��c5��L~�j�e��&G%̰�-�F0�ǁ��ag���H�Ƈ�J"u�#��$�bb��3������ۑ��f����`ͲD0��1�[�MQW����}�;��!�j�΋���C�礪�>��l�X���M<���$Ϯ��ڨ��� �j^��9��ڔ�~t�OΊ�r�W�f���l�r�ӯ���$�]b��� U��,�s>�ݺ�؈�����]GĭU�.� � ��)���y L.h����=�c[�KG�Q��2؊k�EBn�<'����m��T���h�����W\b7���x��8 4+��)�[V�ʯ�Xf�ՎTjV�]G!�3�9tbe��Dl�#w	���]�y�9�S��:^�7ǼeA!�OY�g�U?ԕ�h�b�v�(lLC� h�$0R��c�'&�;��2�l��p�.T��ʜS��^�L��Y����A,�*69�i�0�Y�Bx�q9-�Uc8��u��������㖥E����w���}�� \z:��3�����T�>:��L��_�J�a29��#ۍv5�l!0�@�3�f�k�,�b$�,�<ֈ�,�$g���[PIl�7������>��9Y��}����%���LIp��W�ut�z-��>pm���e���9Z��B��2c�����i�6�,��D���r<������*�c�+��G��F}�M1��j£��E�gѽ�Q��հ���R_�J�������g���)���`�$�mR9����U�`�V�X��8&˿��:+q9�<���͢�C��5�7ʵ��W���Ƶ�D��*' ����GmҺ�E���؜��3�8��]:�	�_ҺO����զ��{yS��`�[�3@F9��76��G}����;��v�<69A��+g^�u��C#��fk������E�X���b���h]��~��7�}h���[{<S��K����J�"p�T�]+ԎS�@(�12�0�;~�!��%w�p>%�FVgٹ����j�$<��.�#��]�K3<�	Va+���j��H/��7Sc��F.��_�y���kX��S�;���#�cJ_�$-��(Q�j�߮����ʜ:�JV�7F�	g�`ס��"�NW�'�$w�4�9��B��Xt�۱z��P4���z� ���� y���6|2�p�z-D��_�4���pc�Cܭ>�+{^��^���D�8�S0d�	�m�׻=XW�&L�SNN��.���ppu3͞fNGD�!ź/��W}n}(9|�k�=΀��1$$RX�j1WG���;Zè��4����_¦��|ӜݕU�4��dZ�$J� �;X��������W�[ōwc	A����]t<��(�M҅ҩ���in����۱�ѕ���jr�S��'��p�6@��#�\C7�B{}E�U��vY�� �MsQ�5�����K���R�����D��&L?�e�j�#��▨]#q�.Q
�	��"(�Ҍ��?Ǐ�<��YB�2k���u�&-����!ͱ4�'��螚`F��My�I����cQ�/�l\v=� Ԕ�����#��D��Nj慬�\g?t3�x�卂9��%�&M��9�����x���~�w 'Q��h���	����l,��oP��7�A��'!4����U���	!z�@�ԩ��f6E�S=Uய�J�_��"2.DT����{ߪ5�Y)j�r�������~�h���6@�eh�V
�D��4�����J�J��]-��ơ/�6E�({����oGo��!�p$�sl~?��ƨ�&$ii��6�˱�Wiޤ#����V$M� �{vۓ0�V�m��@>�2쿮�g�1,���T��{�ҵw�)��əiTC8���ï�HD�~F���l���ؓ��Z7������lp��q ���,X_%�ϔ&���*Q�g}�$�&�G�A��i�k�Uև����	`��qE0�R K�YtqL��g�	�$�Y?3^�l ��x��f\���Y��ƾ��B��<�_y4�<�_����w�7_���0oMO[괢��o�87��ݳ���v�>y3�:�_4�i�J"��*ټ����H�]ltw��ݣ�g�PC�t���k�-D)�j�w��2�\��N��E�=Z��X�P�>	��� �/���a@ɬ����.2�����t ��J���}�A�������9���b�i"Sc�qD|�ˑF�:R��#dq���td$%y"�"Z�kYY%�Hn���Ĵ�OgSMנ�W����RVJ�͓�p���Ên gCi�ru��Uɐ{��y�Ģ�J��֎Rc�A(��E��}���0v?0��U\�KªM�A��<���Ǥj�c�vI�>ɶQ�y�,� 8c��9:�I@]^x��<@%z�C
���q_ر�sTT�#?( ȏ��!'9j��# sE��͟�d[���D^To��K�ı�,Z�f�b�p�{!d�_�h�`|���6�2�c������ӆ��{}�EG̧�=�Y�i�X�d�:�X|��	���e
v���>3`]�!�Y�������A��MA?�*�Ա]�
뼿_a}/�vRo�^�b g�#��!(yZg�k�C��Ӌ��a�"5S9�I���,�\qќ��Q�U6g�8w3��g�eӔ*`����n���"+U���!	n�-����1���/�@" �O��}�`$X6�z���<���N�:y'܃���P�eZX�1 �d�͈�Qi%�7y�\w[�^��y� ;S,,���#��#��n��D;}���кlۊWv�6p�K���:D��t������� ���p�ɹȔ&Stfm����@]��ͬ-*ĸ�t0�6�{F��`m��l�Y���3)%��pB�����MY�;{T�O��;34E����)��|�K  'z,/�v���M���x��/[�u���=��}$����~������b^1�n�H��Ȃ!�ԫMy������V{ř^��PG>I��O�S��������`���e�2�0�ȳ� �è�3KD|��O�d��-�BK����������K��kh�t�W镚�d 1#��6�|��(!!��u�<-�tj�	���Ry��<�lj�a-�m%��)墛���S���f��P@���P�4�|�|��kd�Oi���
� !�Z�V0#^���:6��r�h���y��Y[zO�x5z���k	��vţېywV�"w��C��)�*4���{�7�D�N�M��;�s�lI���7���8�}�aN�|�2g
�/���
u2�a��m�	�>�� ̹��!p�P����%��Y���ajg���B./A)ӄA���J'ݫ���dTwg���Q��Y��D�>oX��.�#:��T��[��zҵ�ĸ\t��d���ҏL�;!��A��y��a�m�$�x�l�%��3!Yp{s:J>5����+�Uخ���I�0N��hT<>�QE]3u�'�}��G�PCaMn���i��m��v_` �$V��?�t��$G����6IpLˊ�������:�>�7�[usJ��9��9�NTh|2O�W|1��}2gB�A����煒������ɘ��!�R�r���W���Dd���0?_&�Դb�
����h|��t庰�Mei^���
ŧ�
��8��+	��,�k�}�,&�]?=L�h�L�R��a����Ƞ�,��ί~#�_�L���[�^��q��с`#�r(���l����")�%�ke��Y,܃� �g�x*��X`��c�_[�G@w��"��L����1ֲ��#�T\�Ϸ;���	t�w�>��^q���K���b_�V�d�6��M�g<sלK���|�������(��p��4"� p�>�k�Z8��0F��4������ ^z�<�j�ݔ�Y������`k�*	�?�����)q��3d=<�%7��k�D�����X+� x����&��o*���@�+WJ�G��Z��a��`�H�^���Mh�8��H��L��`9范�X��%�&��./���]��PY|�:68�5�T�OFt���b6�����eú�_�'㤭��#�m߭���$�e��89�5��Y�	���KW�.2ʢ �Ц9��"Z�6*o��h3͢f%۸2�`y:��~̣ą�8�?GLZ�������/�(P���������`4!�iwޮcRf�=)��US5���f/*Z�:� �N6j�K|�5�m����<��$c��	bw̼��D26M_^�>��ˠE��)Ω���-�6��ک}׏��,�P�%S���,��&x�����>�*���J��J��o`����u����e��Ҭ�*��D/ 3G=����K=�zt��c$Q$^�d��T�����kt�~���kq���,�x�<q�p�uh&S���H�.Y<����̦TMAv\C�se�WB-�Һ��es6�|�t:�k�<��gmi����ӏkJ]ԾS�p+L} ?d>�A��5�7�Ě�5tŸ�x���[��4?�5���DC��S`�=�^����=��z�N�5r���"g�?��A�86��f���܀���s�������,�]a������"�7�����A�c�=�^6,C)`��S�C9�+�v�U���|M�S_^%�"��0C��<[\����8N�I��iۥ�mx�$���*������G�u�f�T��Փ5*t H��%���a�ku����9\:�b��z��  ��Vz?�gC�@�u6�+҈��_�ɶ�W9c锏k|�I�r��4�m:S��5�~6��{/y,�zRR���X���`|2\���vi.y���u�P��Z>fKC��~�#rā�]	y�7����$|w��2'c2|כ��=�:����,#U��
~Q.�H���j�a�&�O�I�@LK������ZT�99+7�b�	 ���;\`�d�YW�4g=��������d�!N�,]�[���~vY__3���;-�����IL�u8�= �����Zڦҟ�M�T�#%vG�hOӃs.or�P���0E��	+��8.]���;�tg3n`�X.��D�+EC¡�2`L�B9��c��lvr ʵk3�@��m����N��N'���q�� �t6R�F�;>,�	�'�m���\6�>��pX��.��A�,Wd��WP�<��� S(	�i�A�A7�yjF2){�:B.R�ŋ��Ǟ�k�"g�n�Q"T����[=z��vs������^���d���A��\��lJ��J��
6e��M�}���o���cC�e��F�XT&�����V@���z�!�H�7DǈJ�t�.�w�`WY'��T����"�M_#�xue?�[�z���O�� ��ds�cA!���T�9��,]�>�Y��~������� ����������w�4�����n��V&�xg;�B�̢��[�J���_P&�R���U��∩\ឝ��c&��F�9�@Q�������Ž%J�!P3���).���>.�U�g,�J�G~E;�Y��_5��.`�r�ɛ�,
4S��j�BC"���MA7K^[��J����ߦ���LTj(�v�{��=����f���q {��������j	�mʯo94i|46w������妷�V�L���T���uwz�ȉ�f��<m��(&p$�\�^ᶍ �W�-ܳ$Zƹ�V��eÏ���T�K�,�Ln�(�S�:�J�Z��eO�^Z�s���D�1o+�"�݇��AL�?��xH���}K�V��G���ԆS_kT(����_{�z�~��,UVg�>Ł�4�B>E�+@�nfS6|�bq��y�L�;����Ǵ���G��ǄDB��ᖴ��nQi$:Q�MA�/�Al�uo>�˝��
 ����vB�2݅P�2\��Nr"���T{�h��v�;n�(ܢ=7i�-�<A��d��X�x�pؕ�߱�Ic>��g���J��f��yi�E+ ��F�G�T��N�w-u@���Ve�R�)iG�s��uz�P�3R����:��u�S�&�[�}�	r�/�ZXU��)��a��A�B��	������Ψ�ep�&+��ٱۓ�o��c�	���-'�(K%��wU_��$[8Y�L܍kb,A+�`l7��3C��л�z��� �ΐ�O�t�Z�DN���֖@��xrٚ%��Y���CC�DMهq��B���+1��YhI�U�2�*�����q�U��xC<��x0$3��Dȍ�Y8��I-������%�m����>�Ȣ��-����1�Ĭ~��$��ӄ�d��/�?1k|j���˼T��c�ă��g͕��.ŉ����&ZY�A�z3�
~"Q�����{<5�0zK�ǁ���`���z�bBU�g�\i�Q���h�I�~ok��ORL�)�`�p�����0��������AI�ßA��6���ϕ�DZC���\G+�_��as�~��8���U\�� �^��@wku���a�X�4�2ha�z/��OO{+{h��.��Ȟ�C���d�㪓ei�ʼ�K���`f�,G�61�Db���o��~�ƮTb��}���(v5~��?d0���@:9�m����:�b��O�j�Xx{�a&�1�oǼF�f����+}�	?�H�p6�����ѝ	������5=�%�QgE��prN���hw��kI�"6D�6ކ��j��ގU��0�A����,�*@$��>�|��Q�86G?��na7i���&[&Q�]K�t���'�쏬tt�nY���}��f�_��?J����׺^��V\�w�eP�g1�U?.>�f��b<XRӰ�̟Y�����\�E_Eq2��q�pX�"B����6[1Y��#G���"���P���CMX2Wvï��
p�V3�*�h�}��5��*�� Y��Y�l�W��Z���>�w@kx���qp�]�ܾ3n%�c>�4���VDj����_ FL[h5E��~�R{v�`P�?Է�T�K��.��h�{�0vBxr����� 2� Wަ�mcH��Ɲ� $'\XsGZo�K��:#G^����w$�$2F�J6e�I�v���=�ghA��1�]�̈́Z��C�c�{v�mM�Ozn�������;�c�[��ZXJ�IFݯw��I�w�_2߸�Gx��)�{w܏�6�7.O<g�d��~ˮ��ⴐg?�ҭ�tm9��i3�����޼M��a�0�b y�d�݂hn_v�4�EA,���Í 3ȠWs@�$;��|g�rd��B�x��l,�q�#9#�Mer��Т'�4���6��A�4҅���[��Eʪ�i	-T;��\�t� � �dAaٜ����Tv��ƳvZ�#�n��)��ҩ�1�{�E};�����fJ�F�}Ӆ2�U��a��p�_�iRR[$���{�y�)�f�i�Ų�g��}�!|��މ�ӉO���*5�j��w&�ؖE����G���ZeCJ��7��}��&0i��À����f�n\8�o�.m�a��>���x �b.
���(h.1�n7'5��ކ7��3M��'�"Ԧ��{+���pE���_�P�!`�d����S~����l	]gSB�{���9^X2(ةRi_��O?�q�h�g���ԍ���q�w��آ�JK�zF݋���.У��g���@i�
����M�N�C��'e˪D}㧪u�?�d�sI�*���iݧ�����ɧ��MoL���"+R�����t��"v�{0!�cոyv±�q�j�@�gg�f%�������wY3*j*Wǋk;0�/~|��ˌ��#�!���*B����>TtB$ł\�z��6�P��S/2�Ɍ��(�W�|Od��o��8���Ü�������������~pD��	4����C����e#m@L����2��T�ǤE�� sv�_��gޢ���˫b���oQ���eM�n���z'O��2�����ƐF��׏�T_��bװ.l`�e
�-7u�>Jbݡ@h:�ؘ{׹`+����S��j֋��PFw�����d�J/����1���z~��;.�J#���q��Ŕ%�����k�ф������?� V^hֆD�=IO��4(*��Hc"Qޡ�3n� ش�5���|g�$g�oh���=���_+�T�8!���QO=_EW~�;-�6�=�]�d���*z���0���e)��:z��.r���!������C�.l7����-�j��2X2��tg�!E���A�o�e#%�cy����G��K+�-#I���,{p��#��Np=۝��i�Ĭ9Co]��HgD��P���֖���^�0O�7�aA��na�WoWr��r1䧻������x�#[[��;��Hk�U�IFAz�w<��}2]��4�����T������+�oEF.5���8�3^ݠ�5T�&j:-p4�W:bsr
�����Y~B0˜��� Ii��6�֡�v�tp��]Ag!�4�Ҥ��o���uL���=���KU(���jga�V#�n�V�MvE�}x�6��Vv�I�r2���{ �@%H]��BU�@��A{�P!ٮ��	��>I �°���nf��lrSq���NWu��`��ԝ�]�#H>C@k�˵�|�!�$;�*~���o�x�w�%]/\��0F������i!X,�cQW=֭Y��%横%��[���]�6����Z�W�t$I�z����p:X��hS�rS'�N �Q����Y4�"�+���C���uG�j��_��3,�Q��Ld�koU�x/��7��2?��'#�� !� �J+�dy�?6�C����eQ���)��/I��Լڡȁ�R>Ŀ'�+D��R�����%����~�p�Xꋅ�Ek�2{�W?�_@IXn�sۦ�K7���S��Z��~a$��2��Z���>��Qp������A|ρ�=���f�q�lA�R��> ��mu���G�0���O~��!a�jKvS�ZQA�O�TԞ��.եη��?�ڝ;&{�؇<RX��0}�L>x`\��k4\p"�n���*���P���?ھ��U��SR��'�Fd�TRp�]U��k��Ѩc�|��gz� C���-nJ�F���t2��H��I�5gukW�q�PƱ�����m��a��'��m���-�a|��3=j�݀/%5�)��[���i������Yg�^裄9�^���ᝥ:�4�P�yC��D�>LmZ1�/"��4�>4��w����ķv��غ�����|���^Y7�?�d�j���
��I�bz�������1tֳ>�o����J��ȥN`��:)D�3�������w���5�H��miUP~�g f�;�V�u�/U.�$����ɏ��H���ːn�?#	�i������\r��`�7u��>�X/�Q�[K�xk�)ֳ��g����#}`�>a'~@{D��o�a����z2�e��_o�4��d� h���J�k�b��X���a�hUL��n7�)v��s7�����@o�x�H�!�*OB��o�XR<��J}�������n��[t��ԧ\��<��{�L�U�| ��<#������Z����(f��EHSW��G$_�
���r�*-,z�)0�ek3C�<���h���w�ο�
|a���{Lq�z�ay�_����G<�-�]��yo�eO�T,;��s�^f<��֙�&�{�Є����/5[�k�mU�O�t��%�޻�ea?�<	��c%^�n&F�����?� � 3O�B�5�ybQ��L{z=2���b���F+o�݅�9o"�l$��؄������^��]�����������-'bX(抶@ͻ���|L1��\OuկbE��~Ǻ����B
P�T���M��z.Dv%�J� x�=i�mq%�c��E��	�~Y< �n�Z[Le�_m�Ox-���l�B�osm��VI�K1W�þ�(�i]3�&��'vm"?�1��e���u�;3$�]��Ԟ��je�^�z���:��D���&�����{��7�*@:k��v�������L*�c�=?�tӲ�bYSt#�\V��Ď�Xs �m�N]6�Z�gΠ)yx�w�ͧ.�iq��;wx'��E���� X�Ě%.lwKʄ�?�U�����g
�\6� ��"1=#}0�Ru��i�P7������[Uz-?�D�R�nf{����2��	(JzI隆i�L��~�����Z){lO^�N�΋%1^��~m��>�=V�4'\6\N�AO����JB��z;����i���ɰ麘"{��:Q�g������tm����I~��4�W��w�:,���Кo0xeA?���v[��* /���H_9|�����V�d*dbu,N�vX�-�)3�O� ��|�8��`�P�	@+��p6f�A>�Pd���;�����m6to��b�=��xeG,f�Z���.e�gDd�����2����݇&~�����2y��[�
~E�p5Ѐ�t�(o��)_TG�4�YK��H���G<Y�T�C�T���.��-h�$a$ZatO��W��{��+M��Em�k�wG$R�su�/C�M)ԔA0���>����J�>Cg|�g�	�g~�z��ʓD�z4 <;M��l�s�к�-��X�83��3��ξ�kk�� �a���1i,S<�m<E8أ��_�����0��������=�0��0�I�J�<�p�W�eZ��@�KDՎ"��E$tI�@6�}����/l��4;�R'!�'W����`F�i�E����������E��E���!�Nc��h��T��y���N~�RG.���zHO]+$JPz5]P�����I�u��u����s$a������-�EdV3Ü������S1 
��d<�Aw�	id�o	o��t��*6TĻ�6�"i��@�$� ���sHZ�W7<� �����(u�������&US�u�~O��3)�ٺ,��/���(��c��|0��i��(�w�޿���%���ԙ�-vw�T��]�;V��5~��/�Py�VZ4z'U)h�\*q=��n�"���"|��SQ�n�P}F�j�� �.�E9a,�t�2ɼo��bT�-�F�{a�#_;���C�������ïp~�%���3&�T-��
����x<�kmB����8�P��� ��\���S��]Z
�.��2���l�г.��r�D���k���/A��RUG�8k��U�*�&�c'�l/a~'!�~ʏ��!9ȁ7�;�@�2�vEa��*�H)$9p�gק��}�{1FZ�v�iԁ����H�� �S3?��f�x��<�^�� :q�n��	 @0��M���h!t��`�1�Z���EH �/�pm]��[��e�v�N�d�y�C8�o��{��s�C�91hL�������^�i}<+nf�����*{��b�m{���Cf��'ޖM�=��`o�8�lXj�0%�QR"�� 3S���/�����洱���"{�m���5G�&0r��z���ƒK_$"~�JIxl��L�m��M�#t��-�
��� �^�/ڗPN)�͖g��.BW,�}Ad�T4����� Q�M�Mr�H���$���Q;><۔I�9�l�8���2�@"
�Bbq9��f6E%��pQ-�?���h�n�0P���t;0����\~v��v�W	�{r�A,��# yN��v�HJ�+��1JuO��m�G���5|�_�9uI;�P]
O��p�h�	r`S=6�����Ti����Q� �E7���!�ƚ$�T�.�Q�yq�բV�J�o �+2�#��[�d�V��Z%����M��[qn�УZ�YԔd[�H�����mB��o4�w��?I%�=���B�Q�/���:hfL�3���̱\�iAR���⨹J���r�=l�,�bn�6Ԛv*�\6�0�L^2)κ����A�Y�nA�QX�	.�')i+XZ���w^-�z��hK�'���0ek�+��露ẍڜ��߬�C��5�`=���/d����� �]��eM��E i��қ���[tz�s�ݏ���c�㴽|G����7
��`l�w����%]�9ޜW����FF�W��'�O��±B�d��D*�[
��u�/��s�㥳J�����ƪ����h���=]qa�^r! ^1��J��܂X�L���-�l}B-ڄN+��-���ų�C*��jer7Uz)�%�/���C���ЙHRpW������n�𬈴��6 
CMD6l< _��1 ��D�ɄQ:\�f�vJ=���VH���3�0/���+�+���፬:�*jW�v��6���6�)˄���-�`��M�7F[掠���6b��n���`�5| �@����V�O ��	#f����g\����9\E9c�%��n{TT���?��Џ��Xܙ$�߃ִN����0�s��+��0ח�0����J���&���NN��!!���F��B
:��l�����/y��5nO�C�\t��a,Ց�����l�>�������r���I>ȝ���Qy��<L�pPq�{�鎊i*�Z�[���	Ox��Ԗ�b�%�+�����`u���ksyKg���	jl1���-�6xZA��#ޖ6���$�_~�܆�q_FS��F�|����G+�U)���:Jf�M%�c���=2?4T'`�\ P�9+�k����@W�$���E��8��p����z"�/o(���_�clҺS�?I	@"���۴
ehhm�G%���6,�"���DK�� 2��]�*��=�Fd{�X��7��+�ol�q����h�AtJX��B�y�{���nȬn���S�\�[�3�a�n�N���z?�j���dE|T!�[��¢��1ڬ)��İyD0�{�#ó�1�fhs��99wx	�����E����`��#$��s1C:���y�qt���?O�e��[tD:7(���h��^�_R
c�)�݆.Ju�~6�q�ND�?�{K�p	�5VǸ��K�J<�C���!)ꍸ$�>��Aɜ0hKd���^��M���U�!�)��8���q������U��b�����$Vgy�G���4X*8SLYc�->z��4$3��
~���IV�!߭6v狉 ��&��?]�1��6�	{!�LmEk�C���?
�d/�PeZ���r�o�@�Ü_i�`Ia:����X�͉@5�ٜMڍr>�����q�I ;����gk���|��;@1�$"�R����H@�Q����-cv��}L���L~�Gz��Ix�ӧ��=�.#Z�t$Z0E����[9vz������f�����	��I��]��yu�]����n�Ā{d�p�8��^�[�d���l�f�A��Q�R�eq��nۿ!�|K�;cm�:uTV�P�l��KK�(M���N.:'3Ng�l	4�#�I_�D�钡�f_zN���R$�.+Uk����t�ɇ�B�j�/�������=���!��p��ݼ0K>[��#*G��G�ݺ�V!� k@@���A����w@�h"����r�C\��U��2?��r�
W�U��8����O�޶)�!��>[���� �����zb�8lS��MG�{�H�[>���U%���J�eH"�n(jك�`����j���|�5jw8��c��
O�{����f�1.�$��P��H �
|��b%��.�D�?��Ʊux[��7�D~3P'�b����O� ��裋���$׫��֞�I&�v��>:�y��X��� �)7I8��#�e��K����L�U!���¶l[��c��\�yv�U�!��"0�b��J�D���8ʓ����Yo�L��
�20�� ���u��}p+�L�F���m�6c�vz��LH��
�8Ĵ��HF[��2
���1�-��p�nYl>O�Sj�ݿ�i�m�!/x_o���}rꨞ
���HH	��Ю`��1���IU-dv��f��$C��5��/Nhr&s?�T;�+Ku���b��#bQŵ�G'c�Vq��������D��;�u5�]�Z=�h�k����[�e9lQ��?'��	j�4�tR���j�uQ>��B�Zi3�=㗩XrN�Ds�U��dw���{X�?����Y��F��IA٣�&�
q]K�@eW���;�~�K�W�¦=�ů�)�?�B���O�U���"�}�ѱ4ɻ? �1��S�B\�V��kg��z�������F'�-�Bk��!˪��ɧ�����b�7J���lRF	f]���02�b����� ϻW��2U��q��i����C�4tBv�jO"�p�+�-`�j�]e+z���;�Noo�Sr����	a�q��B�
�D�������;� �>n��5�|/�5�ʹ|V���.���e!�!Ec\�[3�B:1�햱�vTF��{�XB�g4���D�F-��rg �{H�`���|�/����XW�,v����:̪]K'����B��N�Թ!Wf�5c���E�r�b���*WR�İ�w�P�� �}H�:'�v��84���·�7�s0*3f��m�����J�w(?u��?�f��Й���:ӹ��G-޽���B�r V��5���#.��Pa��J�K���$�����\v���ܫ��f�N�*,��޺ύ
�_�,ʴ�J��p:��h����S,�ɸ�z_x7���VD���p�=oFFP���^J[e/&(}-��q�J:�Fr�J�!F���ֽ��^��E��/�Ob�tZ�S	<��-�v��]��8�}j����	�bQ�	�[���S$8%`��B+T����/�_�ѕ߮Qu}����01�M�J�+�ӈG�vCaD���*�;�A
�1�Ur��V����o�K�\�^�+5���y����jZz�Tw��ˡ����o�g���P(��_Ӕ�	��Q���O�9�Σ*ڋǢV�\3� ���x�����:(�"}L�sI��ӂ/i�K%%I����kE0a�F�at,��tQf
�)�̐�_�^�$2D�xȉ�}<[���E��&�!:�Z����u�
��Y�D�{��%.
��G�Z�l(��8����)v5U<�MKq�4W�|�hVt����~�� n���{u��*^��V��.���YMO!Xu)�/�u��f׹,C�D�1B01�6�6��̶Y�L�sM�1��y*l���H������7O<�~�I��zΥ\�Ɂ��{!�0���F)b����h��®XjU��T�����O�M��N+���??j�g����K��-�=e��%x~��NJ� c�eN0$���ݟ0�Ǻ��dp��U��'k�8�%v�F�%�MY��-��SN�J��ău2]��)���T�K�N��F�)�H��h�����W�f����k�ub$�u��F��+Z#}�4>❖���E��|�E<ՊŰ�B��!����.�G��[r�����C1n�V���=�q	���IʕJ~zE�Q{��r�� fF_���w�Lan����?Uh+@'�t�NեN4�)н��ā�+h���@!c~;��"�)K�#�����
����RR6G��-�
|e���&bn�F�!�B�xD
�<mI�u~M�=2y�r2��}�a)x2�GF�8'�;��_�\�:[�ײ��i �ȑ������mA�yp��
�[�5�_b����i�-�},\y�@q@wr�=	y��a����4����n��И@�i���F.��4@�K??��j3�ƹ����~e������R�{S�f�X���w���뀽[/l��I=&����W��(����YZM���Uw '��E����)�S���DE��2ށ8<�&;:�A��f,@:���U�~�� ����xhS���� ��T�뷜��Y]��a�ʆ˙���3�">����y٦��x���������x	�`= �)�pf��Z�Κ�[X'��T�����G����:B��C��Ss*�!:I�˳�!N\���E�m凸}���k���$��@�E�CwQM���t�+Ê�6=����r��p�)c@�l��HV(��/E��_0-+b���=~(�+�� `�3�B(m ���չV�Ivd���wF���^֝_;ԉK��PKГ QI�Q��%�����Z�k-�	�����b����V���g7��V��n)GC�F��ޕx��y�B�P�0���t	G�r��j#�˗gJM6m5� ^�����I�b�r���4_ƫ@��j��xM�T�="a�Bt���!�
`��)�N�_�Yرɩ򜊒>��%��:/�$G҂j��Q�`J�1��c��-X��b��}�S�oV��}�h}{ft`�`×㘘lcD�rm�r��9��}��=]W��
���I���|T�=�2��ł���*$ygi����kZO�����"��f�t��Q�lg��d�r�X�X򭠽�?�!]��7ƭ5?Ⴀ�[�{i���	�:��;�%:�buSgR���c�n!k���k(��t/S8��{��c��s��ʎ�I@����y�6�nq�L���a�Q��Z�m�p��*@��Ջ��Ϡe��B��D)��Z/�����߰�2�F-�8\�ڙv�\�~�t���Wl`u<�	4k�:.�`_M��5J	҇5� i����[uq���������@���9m��z`�,<���!�ѭ��D}.f{�yv�� 1(�.�ꛮ�O�%��@{�3�Q�'%$�	���s�h�wc�A�Ѣѡ@n:.�[r	��ܔv������_�D��^��E�sVs^����V�<��B<�7���7��8������i���@���W�-��s�I��yG,tC8�S<�5�g�k׮逖/Ѓ�#ƍ���(:�S���MY���6\�=��>��[��I�ڷ�L㤡G�<�R'�����AN�,��9���p��{ъ���/�(�@��g�K2���It�����׎1���MH�p���t��2�9�O(�d��A\��t_��BzTu��2{�S�P�y:=�JH����f��V1��`.CP�% �U���R��s�n�1�+����M�r��ƕ$F�5g��?1���Z�;$�IJ>i�(zpLx�~����vg��CP挑Tg������8?� �йvKX�]�}�A����7(���Gk�T�����vd�F�&��f)��M���;���i��'��%>.���v�e�z��9���d�����%�H��ɍ�݁,�$�n�A�ʙ2�1���t����-	��ȷj�HE��fGCy-D���D1k���|]5]:��oJ�ɥ�����9�.dB�������p��`q�AIe'��7�s8�t�K�������d�Mb�I>XB���^�h~���<uh`��:X����0��_�(�������[9���`~�����˟y_��s�*r��]$2q��,�`j����loGo!C��dT��"��El�E�x�%��8��+�4�����J?��Y�+l�}���!{՜b��}xi��U��x[S��Nl�G35��̩�Ȫ�n�N��x�7.%����}K��Q:^g�pS����䍡If-���UuP�x���B���C|�ļ�����M���ε�HB��0�{F��=�<UO��l�	�B��>aj�X�M��Ke`�8��8o�t�^o�_ ���]�b�^���~�xw62�ei٪A/ͨ ��Q�����Z	�l�b�x�x�#ʂ�������"��|�D���������>*���-Av=�~�&�b�nɈM�ILҡ�ݐD�d���q�;�A J��� q\��X;77����v�c�F�M$wf������ne�su��5�庒��8���)��\��OH`ͅ)���=�O��Ix$%�����ZE}�T�K�~��7�"U6{�a��;�i̕M0��5$=��߸W��6��>�<�{��S��dɤ�Y��?�Գb1�JJ�Ygg��B�m(Hq������blQ.("}���(�:jN	�j"����U� *쪉�P\O�2v^jD���W��Y���T%f���B�\rK
�WNx���1��8l�9ioZ3:�pDC��g�T*����_~��YW�g��6O'��kGR���j�7v� |-Z�5�gx��W�����%ը�C2��u���k��M���Nɷ���/��+���Ҡ��N�}*pw�Y��1H'K��(j��Z�]�&\�1�{'����m��g�g��b]�.��s:����XM_+�u}��H�9 �lB��[�8�<JC��;����[�az� ��wR6�H�C��a���ݴfƧn��nV�-2��{���xM2�$H�[���R�M��I,IP��)��w�/���T���G@O�����B�������n���Ҳ[ ENĄ]���plE�����Kݹ:6K�a��3�ǉc?\�����^ ���*��{�M�ŋc"M�^/�,m��<����Y N�R�S�N&,�Ni�Fi��F�h�?tU�@���c�8a�Y���S���0�j����b"`�m	����wQv�x���0��wg�� �����^�;\%2z��h�[\#��Y���o����+�<hR& ��[�Z���ϙ���-w �x�h	�����$]����-(w��*a�e�K�2d��I\tPś��ţP����_�ih�:å���✁���#���X=_�������~%��ЧS"_�vՓ��L���%6�Bƅ��iY~:�0���r�(��j����`�rm�G~Q7u&MS�C�x%����'�����t/(��x�i5�)❚�^��jo��;t0Z�ZM�@c�-g��Du]���0�3�G@�<u��7��{�'zP����(�=˰"�st'c�<�� �5��d�To/�ި$^L;�[�ef�+�}�Uit�k�2,\�	ؒ��~�$2ׇ��=\�v�e!�e���w�l�_C;�(��L4k}��{?�=�����[Gd�-����ZX�b�.4u>&h�g%W���g &p=P�T�9d�����/��v	�Ql���b`8#���4̵8�2�_�6K5���(^�F�{e8��k.��
�5�G���Ӑ�a�MP���E�l�/����9KV� �\{�sX:��r���	O���5&�f<rh[W�Nb~��3(������?4h�S�OSx���ċ�3��<H�s��i`T�S[����ʼ���A��5ۚ����7gE  @<�&�G�1��؇����^4��1�(�yT����Ʈ�I���N7���:�������ݳ�9OV�Ѹ�����A��^�҂]�8�� #U���ԡ����Ͷ7^�ҊD�D�Zr3guiX��U����-
�����D��.���� umae�#ݪ6��`Y[z���yy�"_�b�?��/M���W)9��uO[�^�>K����`%
 � ��@�&^b����|��|���f�67;�ͺ��?�"�Ť�Nα�I���2��#�m��|vW�X$���M3@��U���Y��]��O�**�S�L�*��Δy6[�bdoyB=B!j�`-O�_���5:�_U^4�f�����e��I�~k+N�*�bs&��|��"c��>K�9^&db�0Ѭ�V��׽q^^�}bߵi��~yD�L�_��fؑ�uX�O,Jҵ��2�8̀2���`_c�9�?�����?Nc��[��>U��(�	�#��z3���3�vѠ)*R�C���"���_��O(�л	|R�Ϡ�:��g���Pu[mu���I.ɬ"�)��� �^2�d����(��hAsER��{��t�� mz)G�*���^;�-��T�()���R��@�%W����_�C��1 ��ӟ2W��tm�ÛUC�	`v���=8Very�0C�yk��۵
YȎ��:F�����y�N�k:�m�yT�A��󓗚2�`�-�\g�@	ʝ��;�ʠ�������T0'�pxDʝM�Ia�Y��[Y������]��0�,�h����c_��P 3GWD5U�L�F�^g�7"�����K\�%�S�Ⳇ��8#B3�\�SP��_���L}QO�V=�r��aI�`��~?4����iCkC�T7�$��Kķ������鴛@��6��bI�5��\nn<��� ��Z��ŉ�U|�dN�Fƀ8&W�p�>����Vۣ�d��O�����1�B�Q�;�@�{�o�I�ȳ�>L�ob$�Q��8�YR��h`*�����_��Xm�X��6��\5թt��$;���%y��ȉz�4��"4g�T�q���^�Q��S���Y�C��%���L�� �H8its(I"~�L8�;�[?�����S��� �t��*���x0B!�d{�?ɋ:	(���hu�o���R��mՎG�-���|�B��D\k��	�Gƌ��0�Ҭ��}^� ��� 3�RΟ˸�<�؏�VĚ�fT��+�&�;{r�V8@1S�R߿���)5�U�i�K�$��uI��R�L�v����13IF�<:�yt�3k���#,3CĚ��{� K�L�i�7����i�ݐ�݂��4x�T��s����~}-��7�� hO�x��O�FM��]]�o��ʢ���0����{"�{�!T~/�[Eth�v>��]�#�!Q=�	�r��eLy]s�Pf4��?m��M������$��M�F�}k����%��5z��\m��b4c̋��|�`i����F��sηT����ύ�ڛ20GX�
$�?��`P(a|��z{H߿E�T�`�ߏ��Z��X�`���j2��N�*���*�eX��Y�y
�)�&t���+�AH4h�:��'7{���]��e4#x�����۾��q~!��$˷�� ����E@�h�ǧU�n�խ2�T_��n� =��p�7�����>l�^&�)H �J�8���JEX��[�J�w����r� �%9�b]� �˹{GD;2�F.deϣ*`���7��q(y�|����5���S)~1q����i�����hW=�,JŹ��2>���� q�I�PA���~�ճ�R�J(FIs4H'�Й�pݿ��o�q����F�@;�����F}B���� Ԏ���J=TN�yۧAHɨlԛ|�>zs1E:�B�kP��*q��30�wz�~�L�J:t�ϣ�HCJƑh��&<�`��9DA���*8��0��G\�/`��81M��6��I��֬��ONռU� c�� ����ǘZ��R�~��0����tvy�c+w@���`6K�WO`M�PK֭�87e���$(U�2���.��ڿ��Gْ����ϸ�����E���J[:�Ͷ���H])�K�|D��)��l����.�&��Q����W��Y����`��q�%�{Dt�v��uʣ��q��P�]y�ƫ|��=�!���Q��e�d��8��K6]R)���	�Ҏ�^Ok�ln��;X�Q����r
R�%i>!:m6�<6�'T9�&emD>��'¶3��φ���&�4��/FA=;�:��ѷL<i}[G(�)֏��[^�pJܛP�%����' ��P��}+�t	\��8����s���<���us�\�u��d���JV��B�iW�oİL�d�Rc-�����G�TZ$ݍ���,zB&��L[�Jۋ+���jw}
��V����$|){��4٦�|�!2�c&7ɨ�OlDoz؏��H�ɴ��R�9,�<�G��V��,�)�I�pTyLkK�k�xY�+�� y��_322l��k��9��S�HHa���?��~��$��$:AcӀ��Ij�\A3]�p�����;erJja\���9��([+������%T�`���H������	m믭�Z��J�_�?+�P���v��Brn C��/�����H����і�8�/XlD�PZ^d�~K3	�Bx/��ʊP�U�Y��RD}^ߪ�����P�+����cO��A��ּ;�Q��1�j��[y j�' 6�gWoj�+��qֳލs�Q����<�V�*�Kv% �m=u"miePd�}-'dѳ��Z�چi�9qHԫ-Ɂ�X6��=���Ι��4�D&�֘&��$��i9}�%�J��H�����;e���NfJ�@�U 7O��v��bu�� ��I)����N?�S&�7�@����0"<�ɮ�������uC8N����}�;4�� zӜ��gP�0"WY2y0Mj�JV���`���ʠ�HCQ�gw�0����s����1&�m���.cc{)e��񿜕rH��|�~=���Q���Q�S��EL w�՛U/cJ$���# ��Ru�R�^��O���5aN�cc9�>@����Ҟ�D�S}؃bB��]�#�n�aؾqK�xйE�2]2��~PQ�����\���vY�Gq�����@�1e���k�J�e�m�<�Lt�#s�#D�o�q��oMuŧ%eD&��l��>�W�h�Ȇ(R�ͳ�8^�,IA��5��Ȓ���e��5�]�O��#�3��#ó��l�]��|�K4 �o���y����}r`���Hb�ؾ�b�.&��We���P� 1NeT��"��h�[ڳ�Y�t˕�)9/����"��-R֠Z��q�''O�r��{R�&�Ʌ�b�2��[}�������3�V��RԌ� k���졻������S�\�~����x!�V�Lc�A��߿I��B-�x��tD��#<3����u.�#U�w�G+�h+7�6��	�J��-�;�3A57�e�-�:j�܌�б�W��Y"���$q�p%��B�_�(�T �.]�{[�����x�o�`*(��}��?�z��`���7rS^�-+jغZ����{>��U��xŃ��p�I�\�a�Ą55L���-�i���|���w�9}}�3����j\���w�������Ĩ�f�o+̰�H^ ���l�j2F2̲hOq ��>���g(鈇��-�Ps\��;^�(����
#V�#1�;���������t��B��`
wi�� w��'�AU�����3�P�p�f	���H�Q���es��Zw��t鐃��y=GO��f��RQO8�6�����&Qw�������P�b�MJ�:2P�w"�^A"C���A�##��S�3��+�{V�D�he�L�H)���R�<�b�9F~���4L[?���9(9^d Ǯs���]�އ�;J;´l_��EN��:��RV����K���1S��v�9@|*��Ȱ�V��q�� )��b O.t+��uEȻޟ� �C$��Gf����X�������䑰W�D�#��C�T�U&�la��}��N���n�1�Th�=H?�/��L�^(ƨ1aȱ>���uI+�u7��]�6��6q�����EnzеR��|e6Л�����`v������ˌZ ������V�g17]u�C.����J���+��9�h��NYц~� |�E.�1�9ŋ��mL����&��+�`���P��.!ٗg��-�W:��&��$�fe�'~��ߨV�����R���G��#V�71���t&����L�r���JN~"xt���$��˷MIѤF��c�!7�մƮ.{���yjf���(D�32��1X�ja��͌[���SA���Գ���uM�wh�Z�%T5��(&��jݓI�q9����OZ����>;��LX����"Q������~���y 	�?��3�2^�iT���n�L�E 8�S�2(̈�*a� r3�M^�tZNbO�P�G�Qg�q~+�Λ]�jQH�6��;��w�NL8�1ܣ��WՏ�Uy(�����H����d��%kJ���l��Q�F6�K�<קV����)�>:��y����f(���{�zؼ%�Q0�O�&�Ѧ���ua�OjBQ�̗/���}�rub�����j	Z�Sc��U�����)�=,�}~�`s�;���{�K�]K�?�
�q���{L����HeHu��Mp��%)�
�-i��)DI�iM��Vc��z[���Vaa2dp!SuZ������(A��7\�.̀<�s�q��б�WB���$x�� ���=�6t!u�_��ZJ�}��`��9`\�Ѿs]��_���.�*��@�c�ܘ��3(7=y��7��Ԋ�<r�Ŵ��#�jcE�� �Zz��C}F�[�.t��+�y&�a�?v��'ۧ�=����:�i���	�)�m�i��{jY��~�����9� n0�{���K�2�򩆧4k�7���	Y�ð� �4�2�ϰ�2�A����'����L
Q=E�G�!K>6j��nX5��[�O	�V�`���r;|��}KT@t��m����(��h�'�y��)�J#[��/�V�<(� =�PRe����6�X�C�F�%O;���F촠}�2�wm��IU�<���K~^�"����OI镧.[�Х�#���k &'�K�j˃�j���ɥ��t==a��'��&N �x���R%0x�Z_�=����59V����w�۝�k��!08�!\�<����k��Z�a���4�?0�<����7N�y���:�!��"�A�|P�Y�eҭ�z颞�Eg�/��6����^�bsevq�4��u]����
�0xk��Qٗw�F��{�5�c;~%u��<�׹v���X�ypY��:�G2gd� W^��,I���#���v#|Ic�ָ�b���%�{U�S��9Q�E�q3*�7rl<(���?����>n�H^��%�1��W��ϴ!dd�$I�e�6cЛ"��>�w%U���M��B�\��q���w���E1�(7�n�I��`ù�Hl��&@���3^�F��=<�կ����B�&��O�N70@�/�gM�a L�j]�����x!�������~U<5s|Z�8�9�0��Ώ�	�� ��V_�����L��b#k�_��`����wX�����3e�U�����svE��[�?^ݻ 0�4c\ަg��M	��	K��/�Ƒ���L�7�6-���Yp�]=G-���z���,�n:*Wֵ�U�N���G)	�%�Ff��=	��L�`]|k�Ɛ`vtu
IL���U�>��a��'k��fU�dB�O�����s���5-��=����E��svkSw}����b�\&�MD� $�����o���A��a�T�ΡV� �8½#i���dI��P�W;�u�'4~=Ku�0�C���<h\�6��-�:������4��S�ɱe�8O�ƷjFfFQ�c�U��M!��n��~���0 9�^��(R�uÀa�i�mȦX_\}~x�z�*٢.#�Ļ�l D���側)0�h�X���z}��s�6,w���Cǵ	��v�
X��p��3%
���[>~)ˍ������4e망x0�vE��tη�|��_T6R0X�r9�U�����j��X���>
��>�2!�V�:z3�wM��D����F�;��@�Pp^��JWҏ���ũ�&�ۗ�\�J�##��D�MḨF�3��������w7r��+���9+@��x����᜖	͗f5.�]oS���=�if3K��Hc3���h��j�����o� ����v�?����|��)Ѻ����ǖi�Gҭwx"MH�v���)��N�@���
�� ��.���m^~�l�!8D�*C<�+�#v��}��F��M$����h�D\����
/��D��.�;Ak)hx�G�aI�ƭ�c������=�T9~EeB�01 ��'B��l/ԨbjP�i�BgHq�����E\�:��J��s:��&&@r	������{y�v��._^�g��Pk[��3Ē�*Dx�)G0��b&�g3���N��}V1fr�E����n���]���M^�Q[�kK ɖ�嫰��s���= �	����.�R�$j4�<o��Ո���H>�� D��2�&���p�{�T|y�7��"P�z�\��a��{]��	c��5���@�����e�e�/	�2�U{��v���&�XG�rjy��Q�9�H�����O/=e�(�>�v��W�yM��_W^_Q�� K]�J�<P���� �P�Q���ޒ�v���cqÆ4�^K��|��D0~U�\W��n���z���`)$T�Ж�j��2(�-FA҉���W`��/G���\�r�c>����g�*"|�;;$�)zP��c��TL-)��`53ƣ}�,F4,�%���v�jD՜-�[h����>�����0�����!�|]!�3����& )w���~E�Go����A�D�;lahζ
�0L�}}\c)�L��o���~HH����n-�A2�����KqFR%��e>A�Ц�>E���jB��s�{'�H��0M�����r@)�A�
l\�紖e��:��4&ĥ$�bi��	����Ho�T��*��b�e�V�t]>S^	I�K����Ҽ�q�,����Q���+�|�Z_���H�S|M���@ )�@�R��J=(�`��ǿÅX)�x�$^#8GMO$�$Gܐ��{bR7׀��(�/er  ��^kI:�V�p����z"X��a�Siߕ�8�t��mɕM����U������Dya���	���m����-�9��l9���V(趋D��G���I���|)��Ǡ��sZ���ةu'������p�bF�䷳����g��Ŗꚝy��Dyi6����_zV��씨WS�W��*K�{�N]��2Ku/���I���)����TK��}��n�6�ItطM��($+�@3^r���x�lZV;��͝�=�gQ̷�� �6��@�$~p'y����\T��Ч�n%<�%���m;q���1��ᢡEQk
��z����0�A}�B���1�E.�[^������|�c׫�V�DΩ��"�^��&?�g.�VD׺k����c뀣|����	(9����]y#���,*T&�����&͖��7\�D�����L���!L�h�RP-6e��Ĝ��/R��e�Q�&N�)^UO�q�j���e�C�q9K�Y���p�ǲ��x����*�mʳ�����jYotZ���A�u�������:� ���Fݺ����^Az�r��3���T�ރ�r(SFɍ�2�?���Ug�qxf��ٶ<\�#"�����AT]ExeT�\4��_��r�>P�Rh�f�ev����l�onFO9}u}�)���ȭ���gAD�)��I#��I2{%*��pg�wl̳���Bܮ��ֺ�������"���r�^T:˴�,�����8�SVk������������d���䓋�5��¿��Tј<.鵗R��]9��;qV��ЮP���m���/�d��$��w�v�Z���v;h���Q��ժ8RO�}#��b��Bl��;*�M�9�I{�q��'e��%�� �v@dﾴ���[\v����6���K�J��A1�=�n��?i:ۙ�V�h�$����������c�+��O�)�N��d�r�<���XQ��D0y���D�)�f�Bb������sJʅ�|~:�bq�����.<��<���(k�mjܺ�y!��!�M�X :I͓�(~B
��Hg��
_�>Z��+��ue�#O?)���AE`�|%Y&Ԗ��;���v�a'�S�Ed0�1 ��U�p�(�*'�x���*g���N��ؚ�|:���R�\�D�";9��� *e��#k3TŦ�����A�Ⱥ6��isf��a�\\�Ѐ�I�$ �Uҷ5���U�;id�$����Z�/*��Ԉ� ٧�S�����P��T�	J�l��Y~�����`$�7��N��+Q���-%�L�R�/�1��-�YrQY*�q������7�k�d���Uf.&+�K!�2j/� ��'=�L����%y?�J�M�B��WО�謩���4��jM��1;Ġq[�����T��?=L�f���{�m�+( ���cv�v҈雩�tZ��I<��^�(�}�#\(F:�}-���1�����;����ݠT�9B���5Z�"�^�e,N6���&Q7|�g/F5w�r|�v�OT�8��>�n�NB:�f|I�7��"�XP��Rt+r�{��*Ӎ0�Vo��M��l2,��Jȧ�cU"�ʞ[�u4.�	j�O���>F���̂�Mc���5\���l����?�1�+u;�8���j�[�8��1���5��~�չ(Yt��q�:$qB$���6�g|�(?�n�WNV�ӬE0�Q�� =4l:�ȉ��)�R��_�Y_B���3�K|��i�Ι[���4�s�*`4�����햮���i�5��'+:E��O7A� �ٟbÅE�L��"�3_�z����2j�P�'��2�1v�Ph��[2�b�9 ;�(cB�|YC_h�*餜1}N�����Ѓ�K)�"� +�l�. �ə�hu������9��{{T
nא�eě0=z���{Gv��q3��4�(�<�ᇐ�U4 �^�K�Ϊ��$��4�B$�����}?3�z7HoT���3tF5��/.���C(\c�Q���%�Ni\I܋,��������������~����d���LwV->N̈́�u��L�7�z�;����ԏ�Ɓv�3��d	��g�S?����k�hP.���b	�� �0[���/tJ��c*�˄%�X#�Ű %����$ #5�X8�����s�Rc��H-USɯ&彁���T]م��¨�x����N����K�_��;�IB�_	�k�̛Ό��
�"�p<g�b��ԘA���+�{�~Q�f�@���~Τ���ɳ
00˯܋({�>�����<\ZB=�2}�ڄLŶ������v��PW�T��#��(��S���\�k���I���V����&p-�i��D���0*�� ي�<��t�֍��e��a��ۻ<|}i<{�E��q�IYe|��E��e�l��P��OJR&X�o�����$��9Q���;\������L�?�%����@�*:�%��9�uhK�)��:�c*�Qk$�m�:aI�0�����+��+A�	V��[�_^��3qF�ɥ�n�g׿�!����;* �So�,8���EօLǋ3E�[n�;H {�\l��ν}vV�n.v�p��Pc�	��� �����r&���sb߈'J�_�G*>a0/�����3���b=�p�u�Z�P�4W��Ja�l�@	�heE}�a���R�ܝ�M'�+��7�s�P�o��=���O:��;'��u�cZW�J*�.H�x��/�+��a������p
!F�=���� �`E�2}C�{X�⡊!�ǌ��ظ(|=���?�����Hb��[�P�k'�t5Z[?Y�t�p�"y�1���Ƌ�ۂ�c�Qo��$��/����,�_��_ۓ3X��̀K8�V�?�nj�o=�Dw���H��:OO�� ���Я�A�܂���f�G0a�MN��XO��$�
Ѕ�o5���.[1U3��V��­�]�&�q�Z}\ε�.T�H�}��TsBM�H��� {-���P�e�=Ƣ�@��RT�FF�I�	t�x��J��=�e������i�@C�$^�]�"��|�X�*�
Qb(�xN��)���/� ��=J��~��'�:��f�nP8]7�c[�<��>���i�����}�m����Ѱ�$ߒ�>-o{7�!�~���`Ekq}vg�	̟�HĶɜq;ρ�!`�Y�%�^u�h��F��hZڇ�����TO��
�o�G��>Ǚ1֙~*���-��Z�ء@.t������$R��kr��o�zHE���X���V�Jؒ�������x�kg�{�ւ���)׬�CWOb$t���d" �Oj��|$��E=/u�-b�ՊI���۔c�_�X�����M����y�%�KW	Q�3x{>�Hʄ;��7Bݖ� 2i�x�Msm��\�,�A�g��-&��Q��i����y�|�W?�������l���X+�ZFGO���=�ҽ��ɩ��L*HSX����/)��<�I�p�V4E����d����y~)�����[��??:m@��١��8T�hQL�ǃI�3�l*1K����};-�?��z�>h��ذQ��h�n�^h:57c��$@S:�3AL�K�T5�L��b�m��
��%,D`ҩ-#Oe��ݞ�.����IۖN:e׼��r�NL������B}w�+�UE���dG���V|�d�7�iz�!�ߧ��u��v���h}��nk�b���u��yR��7|Aw^�#h�aW5[[�Y[��<q�w�����Fq���qLA$�~��ǳ)fA����6��9=	�����~ځ� A�L�q��r���c��g�����NLSX��]����{DlI ��`vZ��&ՐQx�͛	~�O���E����"��2��������Ԇxm��@��c����������QQ���	v�-���(�J��k<@��QpM%� �O�����(��I�ߋ���N���E��$�����©ܣÕx��IA��¤�wzWEe.��*S���Q=3u�>
�,���1Q�q�� \2��m����l����� ��hp4j�N���8P�(ˀ?,<ltm��xd׵��?��(��N ��nU2�-pa]֛eA!�-7xh�����mښ��j#5ƞ�G4���٨�G�Ni��f��6υa�y9.#Q��&�UO�VAR�^��Ĭ��nA��d��eiw������mcƻj�]�MC=bf���T*�o�J0f!.ݚ�ٵ�����1�sv?�5ծ!�mޝc�	��5�~��3��,`%ܴ��T�Z{p��j���:�Az�Y�=f��+���O�[����� ZO�ZO��8�\ui�r��S�"�2<e]�!�-i���,�-��,�'�x*�us~�o��W�Hu������{R�b���ؾ6����-���iQ��A�e�ԓ$Pڍ��6ƙ���]�[�P��}�"s����em9Tj� �d������>���4�#�?ϓo�FW�<֕�<�wh����<�45A�%�1�;51'߀(:O�\�%�tG5�&�>��oVW����P�M ��]g�#�  ~�����φTW4����N0�i�EK�9�����YC�rDݖ�B������!�����tub��$�����y���o���v�q��$�aA֏k������l��b�I`�P��W	��9�X��?T�RS�@�D&Z�R�� µ�f�?r#߶`���!�Z����<됍�*��%��Nr��D�d�>f�D�7_��d��m��)���ȹ�(�����V]���d��!sc]�:k���=2��)I��)�v�i�7S�6JӖl�4��[�8��^tNq<vu`Z\����ox��j#ֿ|�*YEIp�4=-T|�`}KL��9	�0E����`��5O�e�b�h OoIaX�h��Ȋ�U�y�:���F�(�Ab`��`t�y��ad���HҤ5Z���_�H�,ݺ��}�K�C��Y�U}η� �m��x�T叐�Z������ҙHq^.�� �}�@m0�Dm�3o�rC����O9�G٢Sn�Z�ޖ(�,-�0|l��	!n�Ž�qz)�\b�[P�s�����=r�h�K��O��R�E��h���la����BH����"eK=��FT"
�f��"�k�x����	�����+��
�\���Bkă�����b��y�4�t�a2�͒���sW8T�<cL�e��Sk@g�@�6�Z�)���r=(Ԗ�-ͨ���Qv4�^偙j����4��>p ��Qp����$���Y56�AZ6���ltsy�
m�8��5/�掾l �K9�*`G�BJ��k������J���?����(�u^s@�t�!����a��I��
?Z�r�=!��D�T���I��60�X}��lm�>����q��(v8>7i��l���mA���S9S��͙2~��q��(�����@m)$�p�Yd���(m�B9�q�`d��/a�/��*&a�=S���;�nG0��G��%��"d����{U��/1��ߨ��P�<��x� ��K�b�-���рmМ�z���7�qCpP��i�b��7_�N���F4o`?��O�����D��ݕb���:��֭݇\ *��Q1�,=��JЍ�B����w/8���|&�ŕ�n��$��^S_�0K���PWJ��T��F�C[A{���' �����-d^NA��B����d���l������%LW.��(��\�d�����]�n\8�>�g�d~�Q��5�ȏ��A�CE �i���f��&���-^����Հ<���"h�J�햎��E�
?Gw�z����D�k���X[+��M�;�n�gY�L��֊�z*��l�I��Ǆ\�~ZK<�!w]��y��؆a_�&�p��6�s�E�4�5���
7ͽ�h��r=A���;�o�pݗ��*��C��֒��g��+z�f4����.`��]Gb����3s��g��)�"2�[N{A�l��}S��jc<��㤥�y���j�"�Ԥ�;���|F2�)�w���!y�4�mI/���j�<���Lo�u�Qna���6J��;�}~W��_���`_j��/�x�_�dh����1I|�f��#!\*�L���Z�Ӏ�jB'
�Q����vC~>��M�������y�:U�ဏz�.��^bْ��-������#ީ�xC1Պ�����0����G+���J�1���й�A
VͻWz"Ĭ�����1n��<̵�c���H�����|�C<���*㹑�R7��.��?�&�躆f�Y"Z
�]��lԊe̜��.��r|�� ���힇mpv�s%�������4�$Z4��M�ʩ`����gl��p��Z�֭��IjET�$s��i!�hk	8�'�!�jĨ8< �^3&T@#�_�׺�U�;���t� �08J�!rs��B��Ͳ4��A��Î5D`�Ϙ�oq<��.4�h��m���lE�|��σ�}�1����$�?�Ȫ��j��\��7O��`�ߐ�I������˕EH��J;'R��:�<Nha�q`(8�#�c�H�sn�ڊ �E;�Gx)��3���wD�Ǘ����F�<b�3%�5]��8�~���K�s���J,f�/����gV>�4��$�淎����F�d�T�����B���SD�$�0�ԨVE�Arn��w��EnB�]�-�*i�����]�錅�1q?M�>��]�+y��o��v^�j���F��
���GGt�q�<saM��_IM���r"���wً�4�m]�J&o�c�]�P���[�<W�k���_��D���uA�|4�6�֖7gQ�����;ʐ�]�{z+K�~�w����Q"U;�\�mi R�xL*��t�a��r�f�W�&���������Z�r;�͕�4���оjLV��ףE�W�)�AG�H<��d��es�i�<�1����T�+����: ���N�!rn��~�9������ �xd�ˊ	R6&�ާU�pr}�je5Ey4ZW.�zg�J�~�*Bmj!��!8'P0��Ɲx��$�"#~z�H��A�y��b���n�BO	�1*[����dg ��QM_"g˧qR���"��1�m۹�����owԑ��lx����w�{�vد��Ʈ|��~�CEXz������ T"��E��>��V�3�DY���£�>���B%��(�G~��ƺHU"*j�b�:-pt�n%�m�i&��w���q�x�R|m|�DtF��ti����/���n��t(�$/���2��GR	n�R��݂[�bλĜ$n��׋߄�oT���4�;V�-�0;=ud�+�R��Z}�դy�2\-��.o���>�������^:Hp�[H�stD�~��j�TL�K�wu�O����#��<S8���ܫ����j��mѱܧM7A!�(��P� �1i�r��D	Nr�R�i^�W(zy��||'~)����B�cdiD0k������]?�c\afb��b?��i꠺>��e&Ʋ��lt7�-2\����,��s~z-� �`��D���r��J�p�2u�^®Y�H��+�Xu@��:�?�9�tέul���M�-@4ז��<���,���be��͑�5�?�N�9ɹ����A��mEX����"�{S6;s��+���-1E>�Ь� `�B|��zT�`�g�o�`(N�F���L�F�%i�t�{���J,�^<k�.��ů�SA�q�X��
(m2�K��y�E����^O:K��c�Zc�:�hT{?��|�~n�m7����c���������\-ر'��`y��H�\g��f�L�K�������[��,j3�^����栔�ny�����d=^�M���D�2�L����p�M�}�_
'?,?jٮ��p:�3�{��B9��
_��t����N���w�T�U�o߅����_bE�(Ȣz�g���7xiZ;!5��Pa+趕���4��2��xm[Cft ި��)^��*Ҳ:T�f_���y	�}4����
��A����:MH�!m(�w� m�a�2͟~��ň<�L��d�h�~�:.�
���_N^�s���2`O���qԜ���f�>�+g��N�dRD�y+[I�:��ݏ=@I`�TY�F��	��m	�[�Ǧ�wt1D��/�ݏ�XӣKΗO �����W�<��S�\�Id H��$XUp�r����yqaW�V�nU��n�7�2�Q �G¿C�|�t4��?=�*Z�P44%�d�J՟�xI|7��zgrUu�����z�'�7$��� ��)��h�<ڴ$q��N+-�Kӎ�N-�֬^�j�3�ӂW#�"��~�-��m��;?B��� /I���"b�s�8��`����î������fd��&^�T�[��m�*��=xo�v��^��}��x3�A���/�kX��1J4�95Z�FR ������*�l���))̲Q��H�cm�V4�`��T|I�>>+��xaڀ,\Xbⷲ�їoضi$�#�̨�W\,O;��
��\,�k�]���[@"�i���4�ڈG�ۓ9��t���^��)�G�{z��Ȭ�0<�������ES��Gk[�֋H�@��?ot��$/t�B��y�%a��2o�>ʨϞ�̀H�X��6��B�>�oI�>8�-�L��I�d
�r���8�PQ!���o��%����h�>����vť��:���NB�ʳ~Vë84.���תDĆ�6�Er��~g�H�gD3���H_�F��`���R *�f�pxɜv��qH�u���KϴM�����
~X�8�E���m�sv��SXW�����4��M!���ߪ"����8�Cy�h�2��]�����Jj�Ĳ%9J�`������<`|'����0q�}m*�y����"3�s_+6��K{PsY��6��;J�����[{�cD۟���4<z��˹ܟ9��-w��Lی(0�Puf7�!#'iͻO<\��:z�g�8q����|XΧ�:j4O��֑S&�!�09��vק׽�|��XiB�C,�t �q���݀6&���V�$/�E[��	�)�-�2 �;�>�W����d���iׂ���?pfJVa^���XI-�{�_i.홆Rx�o����Fȩne$���7W5L�a�߽5n|�^E��]��k}k�G��Bסv��,[��N�i��r�%���i�/����Pq���^�*�hř���q�t`y�!}�%nM�[�~s� ��:��7�wn<��/�jXe�кb�A��Zٮw}H�kf�"1���u�:e���,�^i��+v؏J;�
}�c��[е��$(��2��� v��q~� �m����X{����8"���Ԑ�a��n��gi��n��/9<�נ��4*�睍k̼i��<�J %���J�ya�������\g@%DW��.i�ms;��c�IUMlˎ1�Ihn�2P�G�Ǫ�������ߪc[�BЛ�*E��׃i��Y��5�%�$�c���ݢL�З�bDBmHJM�o�/��f���%>c����M����]�/*$��*�de����O��~	Y�ӟ� ݜ�[ѯ�B�I�2���*F�^��{%-ֈ�U�x�\'��8�/2����@y_����;��Ӵk4����S:��Õ���g}m ��������g�H���.x��h5����T#��6~_�)qu������N
ׇu3��a����?�������%����(�Q����݊<)�'��f�j�x[{���քjV"���xX:����-���X'S����'���[۴1K��9Rn՘�נ�I�B�FM9w��	cg�w��N���p��.ⰶ>�9.i�fk�s�Kk� �(��%F�GOC�L��,	���Ǩ����p�&�V���������z��ha��G�]x(�)=��@�2�m�C�9��F�DF�$�Mm�ޛMz�͈��'�;�KʋXY���(nx4���u��\5n�i��au��s�$AuIx�;�_�H�����e�$�H���`O�����r���;��i ��A�q��:S^w��6�v�����x����HH����x'��PQ�i�O�.W�s��L��Y�]�Z�Y����2Dz��2 ����-�,s�Z	S�/��je�W�/�ػ)���jo��Ɛ�����
�
�BG��>�3ߦH�+� ��U%��?�g'���M�0ψ�
��S��O�>h�\
��� #�ls�P�3��e��L¬��gOsp)�Y��� P�r��w��O^F_�fD�BFb��3��jb�N�Z�Q��O	K�v�i����ﮈ���6�	�v�J��o�l!�.S��;��|�ڤb���3��ǟ�*C�����g�c4E�ׄ^��چ9��-fZ�{��n��Q�=������Ag2�hB���g`�a�E*<�cW�T�q{(7��]{�m���}�S)5�DH���rG!{s�5P�D��ƫ������)�&��2�eCF�v�C�U�g�!+؛��]����5DM{�v�EKC[1s�hYp`;�HTE�B�VT+$�l�U�
N�~b���o�.��C@R�Iݺ2]B�V|�k���븶�r�B�){��N�D��ԕ0_zI5Q�����ѝ�\L\������HȮ��z�f����fٰ��
T��\���?��g�13��!��(�)��`
t�2?�R�@ܜ�UKF)�vZ�7 8����U�5�hw>�\$F�U�u=�o'�{ҟ��> c�U���m`��z�r��I@���1�\5?!Aj^d�-'Bz��O��1m�HsOTD-��W)�L�g����ԑ�(���I���pD�O(��R�l�F��v�"����l����0aԋ#���s�.�71ŭ���C�J�H�C�	.�i#�/S�E��^�ݜ��m�|E���A�B�\$�▁2���`��Bt4|6�'W`���KA���dͱ-�Q]򴠃�in!�`^Ȭ��<$����D�W�!��nkK�\�T����F�<� �z��B8#;hn�N�ks'�ŬI� �ɭt���ndա����F������av���9Q#��Q��:������H+O�k���y�ˑ�Ո���(2��ջ99�O�)s��_/+�@�4XKڀ�hj �wٱ�"�(cߥ8��h��P:`�5t��;-ɛR*5�ܵэ��1 6�5؋.�� ��[j���͞3�T7�&N	;�����Y�{O�@�Mi��2V&OS�k}5W�Kd��͔�~�_K(�uiG���K��"xy|�%�ɘ�E��H�/����. O#���SվYv	�L��Z�m4�g��q���뾁{��|�p����c%^�:�E��(����%-R�r�TZ�����d�J=4ʻ΂�|^A4����]5S��Y���#:���'��&�p �}4�ol��a�Qn�aѤ��Q#m8�n�;	\Cl
q6����T4.�+	�V4n؛�fѼ�5�,{ѣ��_�s�"�U�j#��A�ȹ��BA��?q����0��s�O����/]�(�����.[��?��]��M��'����"�,��%��#��T�Ȅ�(���gqb�rC������H|2�����<Ӂb�-�swI.��>�����U��DՐn`.VGFB>@D��.�bg�f��Á#�Ν�e6��Ҷ��+FI&��A��f��~gI���[��tٞ�=�h�ý=;�H�UEc3G��*=Oj��?�OG��X���I|ݕǣ]���?�۪�Jj�D�����������#5E�pt��ӳNJ�(���7��i�g�0�5��k��@;[ߋ�خk���~�����L��]�FV�߂=i�J��"cU�5��Ѡ��������][�#������y(�kfl��>��Ő>�R����?�����s	 �2����E�N,̻%m�=�ɀ �#�h�&Ǔ�X�Ӿix�	
_��rC��6�2�*'�6����!�Ge���Δgm�C|5X��-��&��/`��_+.��n`\h+7}j�kt�G�촲Xaz�+p]�˝�]d��#f919\ۥ»jO9W��nB����{n�MW\�3��5�K�g�X�V����?���W���U4U���~��@Q8�j$,"�	�|O�?�A1��ӠI�栏;��_~n��v�/�����o~%�������A^鐷�����|���uT�!��J=�`Ar��;<��G.*eX �Ҩ�(�I�;o�-���"-�o��]��K!5����%��ś���Z7�7*O��� �y�� ���.v)�0M�Ne�?{����zCP2:��nQ V��!�>~ĉ�
�u,\{�%���N����]��՜(QJpuZw��6t �B���W���[�!�b\^���zi9�3�+\��xPbX�!����/_q[ <G�;��(`���ϖ��o=jY�a�3G�b�«mlc�sɖ��J��x��
�-�J^�9r�	�m`p18/#��qy�A�������Ѣk
��# �efi|�&\�9͠�����Zy �b�?����,��N�a[|U�BQ�N�r��Ma|v��.<b���/���(ř��ڣDL�N`����m����B�/�ӏ���~IoR�|�Y�w Ų����(f;Y.��Ah� �ſ_� �Ml�X�9U3���h4
��;"U蕏oAE�#�UFB�Kk ���Sﴁ�#�ȼ���	�� e��6�1��j"^�����n�����.�:��h�[�ЉD�P���\.=\�9�c�/*[�������-��ҡ�3?�Z��W��w��x	�6��|3����%�waȼd��������{���e�k)5P�"G�V�.X��)��"k�I�]�0ǅ��]&�Y���6�R#h�p��^��2��ЊX GCP������u�k���/��W����T
�狮?����/+��jL��d�y�9'6U��s7I�z��/�3�k5��_�,��E�
'E��ZVsJ,���e�<�l�t㉲�?�j��$܍;��W'��/@e�9�Xe*G��p�m�Z�������x.����R�ԟ�S��{��9�!"�r~��gV�t{����@k��*V
����������a��!J�;|��#&*����ː>�������#^�M��XN?��k�@^���m��Ī���XZ7EP;�Ӣ� �����.o��B������wq[��_d���|��;Hm��F���@}x�� �>���m�b/��L�*f[��d�U+a���L����?���.������F5(ޯ����K��s�z�8� ��(�3[jnC�d�iW/��7/�g�R� h4�i���$��.��t��]�0�j�����(7�Xw�e��~���� à�?������Ւ�k� �Iϳ��ɒ,���{��Ne�=���[�b�]o0/�-O��Մ,�s�׀W&5��L����{R���<c�@[GC�� Ae���}Wʾ��V��R������RM!�$��^��2��s?*k��M�j��K�A��rU��Wy��6t�/W
r���_7�pԟt��ǡ��D���#�����bΤz�m�o��+���"������֬ �M�<_%�ⲞDT�l2��R%qAG�U%-a��s�QGǯɄyV=�Cm#���-;��3�Vd�ę5���+5J���p$��ֲ@�_-�H�t}q�n2�gC���!�<^�j�g����	�ba�E������S;�!���<��x�X��I��'%d��b��\�`�:a�3=ґ�y���"�փ����)% Y���<��XbwTp�-�w���)��^�&E�l�%tk%A���5;��7�t�2�����э�d����E��7У�"�ޗ<�����%�M�*��<Bg(�[��3@D�L�k\�c4{��&4����(�/@q@�(�D���g�'(�3�܇N�^B��[�wX�+����rΝ����!V�,����R��v'kޓ8�s�D`>�A	�'�K$7��'�y���_!����a�0��.^)��wᑙ X�m�$4~n"!�U��DO����qɣ���GW�i>�w6���W�=�����F����:p6��P�1�0ۗ�ܡ�Jy��������;�H����s��FTXIŠĝ �Cbd@z���UVX����w䨼9"�15�D�b�q[�z��1 1k��Qa�Pqi/�g��%7�K��MM˴�H�O�ͮ�d�w�^�ztb����?noG�Ao�y�4ߏl	�8�OIP��( >,%���m���$
�C�i��Ծ��ѣ�Ϲ���0���[4���}t-�;.���c|��r�ۖ���?����!�&�L��7�̸�~�X�2HG��W+��W���e�B�_g1�mt��-�O��p(]�VS�&K��lM0�x�\��{}�s�|r{���	G�'�6���6�9����΢Itr�X�U_��Q�>r)�(,��՚�}�d���ծ��!�d���+���XIQ����j/��8	b���ޔ e�yAj�I+��3|����;��,���=(5_&��Y�&_^x>;�,���k��֟^&4�4uB��*<i0Ơо����t�pF�08ZHh6�i���ki
���T)���6�w+_Od����\O�Y	����#����P9����)�����Vn�����K(����.<�T
\�M������#w�K����@��Kr�'Kb�L����b2�#�ͽ�.9A;�99dy`��SIi��È1ğ�z��2<��V����V�g	�"���>�ͼ7⺈a�[h�Z�G�����_��N@��$f!���m'� ߍ��2�]��$2�|��cy,?�:S�#z}��8��1��T��x���
;���@Bw����'V�奉_`�O�o��d�f�#�q��X������x9�M`pvM��P�X�5T��7!�'��*�w���2�U*��`F��!�\JZ� 狸V@���"7�
�X��~W&B����O��kz�ڬP򗊔pm��Z�J���ۉ��hKjW��Oc��/Hk���ݖ���9M�(%^:�S�h�W̡e�דC"`�5͔����T�Ә��Ԋ�����ȇ�]������J��Q6�b��;����X�BgwT����TtZ�5�9e���@���ۗFԐ�aҠ��:��]��� ϯit��˔�"� ���5} i��uY�`���l1H��e�}�$5�-���`�='�`���n�E-��O�<T��h��ysUV_�?���]@U���1�����3V.Wl���+6CZ����wW�RGJ�vP�eҤV�#��jO!�|G$!�?(�=���DޥV�ia�o"��G�l}3�����́e��*��n� [b��rn��L1-��7{�Ǿ �I�hw��xS/F����T�֒�'��:��Y@�t�b.�Q,��0��Ά3���ݾ�~�Z�ʖv��uSєX��є�զ�%|�b�?�zbbG�,�օ��ٮ����Ɨ�nF��p����؄8��4�۞U��[��E98�xc���B�v#���ˑL��0NS�B���UP��;�f��x�)����[\�vҭ+�]�*�
���X��rk����M�`ƃ{�����?K�!��Q�h~Y�]�����t�-���*���+喭�p�>SZ|�C}�ߨ�j�B�c���L(�\��n��������b���� ��%�(��h�GκP��f_nyR�������K�U��t:G�R�����c���ʞ���՚b��,��:C
��`�>�z�y��tm��q�]���5��V�ү���1&1�iB=A<���@M(C/]�E�0CN�E��?�l3�ɪ�k=�N~�5b��_b����+���E��Hu1S�L�ga4t5�f��53�����mz�g���$8����{X�ZTw$3�Y�m�Z�����V�Z��vL4Aq�V�*P��B�Oݿ�WGyF޺$��֪3��-�Vԃ�scG:�Y&���ޯ�Q}�r�a�#�$o'�Lw,v���&U��;W��A� G�N��н�f���
�`}<�nN@X2[�x�i_��pj:lۂ=�y*�&�I���i-:$E*�����x}��V�;t~�I����(�oJ9� �x����T�sܡϐ'�W�ψ���y|�؉n�j�qA�v��'�M�N�	Y��i�"�ÇoY��Mؒ{IN��^���DTW���=y��+���Y!B�ؼu��6�zoo���Q��K���E,¡�]�!����5l�;<'"�	������փ���ʣ�g)�LU����L",��K�8����Z�me@���G��F�Z�����`y���N�v�:B�H��d��J��t����ǉ���L{�����Jq������˫}F������\P��@�FfX��d�J�46��}X$�ޣ.�)am��8rx�6�kg�nM2����?C����N��
9`X�~�#I��D�[�kƍ	�G�E�1��6i��"��<_#�8��D��1�����&���żj�� ��a%��g�_Q�|������#���zC]��r��Mkto	� ;p�ט��z��>W��Љә�uu�\_��^�J�C���N�����������6n�T_��T�u�dd�P�5("��~�?c�2�1%��O83�V�FӃO,�^�U����7ժ��$>�*���ix��x7ij�[��q���U��j��S�z'�묍���g�ab�Z�	������m��0nZ���ܵ�k�u�F:Y'��u4
�J���|���N[���t��Y�?�P��v������Mu����|2����/��q=�3�%rH��>0v*������'o4��G�����9x��.�T"��y��tq���돛�JI����ׯ0�,��{˧"������t���Xx�
����7x
���UEM��.:��*��\�N��&v�z�J�Ȭeyo��Q?}�e�~�#xq�,Z�C��Ǹa�N�Ƌ��b�Cp{���,�8ń����6WT�ǐC�TG]5��Lv�r�������	+t��l���ZM.ò�h=0��Eg�4��h��^f�^�M
�� ���s�۹ TG简� �lي�������_�vEO��G�������7P�����q�Uέ[_ɷ	�nk����.�O%��c�*�
����h����X����ێ�y��'��ri�Ϸ���H:�����{xh6�IH�7ɳ��ѻ۫%�_u�i����zEY<s�Rb{f�j!|�h�	��A�_�����D���:��}"4��Q��>�Ǆ��E�b׹D?ɚ�]/&�;�Y�����6=
���XE����	�y�d�/�|s&��>�{�������mێw��h���jt�d�M���F�����,�nv��=&u�	�8�ׯ�T�ja�gГb�a��H���|�ct�	����A���j�b�}r���^i�*.� �a���]�L$��i��a���8e/��x[n��	U���Jm���H��N��ͨ��� M���=z��P��� F�dEv0��LT��}���=i9�Z�3p��l�&j��)7�&\��v�o9;�Z�@N��9B�I䨜^^�tE����5�_Uǁ!��Yn�ѽ��L��N�h1p'pi���<*��7���<4c��&%�Y`���=Gp>C��)ҙ�{�@�A]O�6�V����i�V�D�N���h���fcOeO�n��z=!�H*.�R���>aCΆKx�R�Z�3���|��Q��:�ڗ=�H��_{J���ow)#;3p�+��o�"k�ɱ*����s�R�FlҒj��]��)ģ�_φ�~!������ڗlL���$���<���{bF+��&|f�.�_d�������R�74 6i"5��i����:w+�Ql��E���B���S���{�d��~>�6���v�P#���n�˖6�Xv~�9{$WktAS�z/$w��l^��$my=� ��I��ޯ��q.��y��4�K܄�8�h��-3�KB�|&����ȓ�6�G��c�h	+�zv�k��i�ZR�㍷���.Oj#�5��$m��?X.TL@�f�e�d�@&���2���|]�i���Q6r��J0��SŸ܇�ڙ/ �!��ᯐ�9��cC?<Vp��_}������q�m�{d�	u:l�V��Q�~V�Λ����ܽ����v&m�u�:x�a��*GJrO��S���<LO,i�X�ʛ�V��f�R����رBvn{*��Pe�=r���v�J���\�m�(g�����+�7�$�F�{Q֬	�0���5+�·��S|�;��$.�y~�	Nst�Ʌ��,�@�wC��DT���vR���\��]��uV��d��=p��uԡ�������d�!
I$���<w(,��cx�]���?(6۾�G�4Jfm��Ȝ(��^G�sv�~)�� �*C��܅�q����E��4���^ee'CH�V+����Cs��釾���]�m��y��[n��vY��6��Y%w�|
R�qAM&�A�_��`��j�ai��|Z9���'IY���N\���k^`�~���5m�aX�)c����ȉ�l~���U�z1.�S�è�}h��ݮі���Ⱦ��T��=�Īo���o��f�������F�jF5%᏶VEȅ����wƍ�ҺF9�_��W����ݪ}*f��oKEjf�{�x�r���/b��*X�<T%�w$�=����P�J���|(���%Hrj��;�jr~	0�����!8`y�DZ��kU=|������%��doH!]yaJH��G������~��]̐�</�m1�;ޟ�6���F��1(�&��H˯��IO�&�"�.�C84!�-�o�4�>z�\Z�x>�h�S"+�Q{��eO�V|�Y	�~�;�9�J#*|�饋�����?�0�v���e���q�/?���0�
�B�Ce�!�;�����{*��n��=�@v�B�6��������pw�tΠ���ގ�����Cv�x��,G������@�Y�c��u�D1v�|I���km۶l%c~�BR�2��.@�@���Y�����Q� f��4��DOB�������Q=ʜ�I�͂��16����z� �h��&��\����>��4�G��&�����#�� '�@;]�1����b�:��,�\�?=G�~����?��g�N���,��"��y'��NF��7R��ޓ�)^b&8UҐ���tM�o�����8 2�B������>��q
w f�\Tb�r���$�rՑ�9QnA&��D�q��P����CLr㩒{��s���>���T�©J�A�yTn�¼��e�`z�eq͵�;#QW��B����D�f"�;^OV{Hi$���.MN��b�'r\�f���=J�AG����U	�1��Q-�F�җB�Ի_�w^d�_Z���L���^�y�ې�?���"�/b�Bo�ZE�/��Ի���Ç�;�н"G�m%�{��R�nU�F�sR���Ex5@��ӱ�=���S��Wi�l&��X�"q�O�Ҋ �>O�5A;Ks���g��0��X��A�q%6<�L�zD��cd���C���?��N�����3Ǔ�|#�!gЄ
(fG�~�Ί	�Vɪ���v@�� ��*�7�������j��3��N���v@�	kƭW�#�G�v)K��Vd�]o�p�c�y��[���cq)0S�(s�Xu�~6�C�:D�L� (><���'PnWJ����j��@������16Ƶ����僇P�M��Z�Z
�z�f���)y��g�������]��^��q)��4��x���/=&C����`�Kdj.q��ê07�I��p�ĄKV����~���C�ɪ������?G>���D�3�Yr�������Rk�
�,�/Z(�m��J��yLmhI��������!;��ׯ��� Tb6���1!��f�JǶ����r&�9��K��>㝀����\X����6�E��6����N~�J�Dmӓ˞n��{�FK���=!��̰}S߇Um79GY%�MU�xL�X���g������ڟl�����=�N�����V#V\���J�ϵy��g�Q-��[>w���/j���%�x7��H�i�,�`x ���Fȿck�����w�����~�z��D�-q�\�o���Y�0� b�'x�a�ي_T*��o�s��'��W�D��W2�|":�tr��ك���b$t���Z��D���Fy�ɣ���>�iP ri����όLP��}PД�p`@	�K�8�M�E�Ģ���VE7d�� ���W�r�;�D��ͭ� g-"�$�8��,Q^��O�F�C�ަ��|������I{�/Ö�q�L�q�s���p���jA�9��RԏL�e(mJ���m�]�x��X�!j.~~�w��]|�~|L���V����K�^�Lv��+��r�>J���x����)�pID(��j����mi�UAY!�Uȡ�����t�j��g�W9>ň�'1��4��^�ƌ]�h����)~|B�OB���]굽�!~I�N�OQWs�&���
�2� �	��.@�87n�RV���	�N�"����5�����	�Du��G)v�0�z���>��"E�Ҥ�P�Ü2=4�SLk�7���"�#�!?]����R��yg� [�MiS�у{K�HǊ���B����&X�<D�.��g1���]5�ɖ���:�ͮ�����4�}c�¦	 0��ĉ�M���r�AR���`���ʡ*�@Y�X�����!T��e���Zb�[U�����L�B�/~������oa[�䴩zc>� �:�0���$h]�,Z�!�g�q��j���/�3M@���K�K7��� �@w ��s�p��H�U��7a�x�K|��%!%Pw%���{�[I� �n�ٷ�Ԛ3p����Y!��aO��\��Q���L��-v�����Q=�/���'<��b��k8HC�x�b�t��v���c	Y�M�܉��Ɋ1whԕ ל!$�̀0	��:3��&�3�xoɋsY�e���C=@�"��0Ǝ����Q������c)\�w<��G��iO�	 �;m�H�i@����d��Ӊ!���b��*��0=����1�"^4[�id��*_�2�s��f8Q>U��+�$Ԅ�OC�+�(�K8��A������!ݽ��6���ꃺ��+���^��(��
�.���O��hQ�h��� W�:�м��cF8f�Ո�q\���t�8���n����MO��Rn��w>1Uq�^�z��n4/�#�\}�v�5O�YF�D���G_�lZ�!�o�3O�z)~\��˵@F�1&�Ù��ܵ��8U�6{	$(��H��7/q�1��˹e���e�S�n(A�\�r)RK�H�xH���;��RY<�&TB�2pi&��r+3���C�ӳ��,
��)��u�1���;��B�Kp  �����*(��錯�7��2�Y�/�l j�7<�!YJ˃��:6}����3��tf���y��?��=���|7�2���Go���H��Ն��j��s}��2���SJ�1>.E��r��po��67VN6����ZJ�7��`�5vd�\�̜w� �=� =��Ui�S�Q�Hu�4����t?�6�%�zʫl�Eq�%5�=����c��������i�&"4_cw��\6���ױ��n}o0�|���Qr�Yظ��2�^�,κw\�x"5��ը�g�$�z�N��HѼ�3��11�N�� ��tn,b�]�;��e
z�F�{�k�<�a�"�����(�+�ӕ���ޓ��ʎ.S�V����Z�珝u��6ǭh/�HI!_�6�{�Z�e?X�-8�iW�j��XՅ���TB�rK�S	��`p A[������Q���~�ع<#q���c��j���K��]�B�MDD�m���o$��6���o-/LW8�#e�32U�\,��{hX����ۦ�3��j6O�u<��23}�uo����Ջ��h�N!7��#�\UlZ�X�6�����a�6�v������`4��y���Y�=�_w�L�\�l�#ڥ͉��XF*�\|��7w9w��F�Ư��h/�>�S�2'���=���An�ĸ�蠂�V7q�����U��qԅC�����C-�0���J��)͌����/������g��ܘ�aX!s���׾M�M�ۍ�IP91!����h��i�>�I$*��2����V=��[�PX.�R8F�2�8b]�R#��c޴��y��!$B��߮�|Ù�g����b��[Bb����y]{ŀ~���J��v*�W��/3>���!��Y�PG�E��
����,���:-"�@�y���ȉ��,l3/X��=hf�W��يӦ�[�/Q��g�Ը��'}�4�y�d
z�Z=İ�<�q���7�4d $���b����^P�&�a2�W�ValS|��.uժgIk����YM�?���<c͠��_��T8����2߸Ϝ�]h!�.J��嵠��|?��A���ۓIW�fk`m]�m���~I�Zbt_ �|��"n٬��3u���6*T��1�MB\�c�];Jz�qA�~��к���
teĆP��Q#���L&i�t�},�����W�u���G�w`�B}�"����;x�OB��9���WxMaE;T�tM�A��?T9�� �|�;!�����@zqg��S�Θ��q@�쟠:�Ru�@)�-�*2K�qqي.�c�/��(�E���W
��*��W%�&��N��\T��/�xɎ�`��_�m	��!ԋC�4K��s�Lji�O�.b����W��LY}����B����%��8V��K�� _fb\�}"y j�q�����E��� P&)��D��M��c�7�/���s��H�v:^������>�wΠ����Z�UT� ��Qq��7QO�;`Vځ�,��eQ�;���H[�|I�0�\�Dy#2KA�@�.3��{0$�+/�n%;^��#Z�ޮ�p�FV��aF�~�lY(���E.E���x\ҝ�oT���p��5C���_a�~���I����ڐHd��~�.RSUp��Y��q'Ç�áB�Y<�+B\m|p�Q*Z�yL���Ŋ��@�2�UOs�y$F�[��i���!)�W���Cg�MW��֜�����`!q*�9dލ?����pMS锺��rHF��Jpn#S(Z��m��M�58�ܳa�j�?(6b��:AdY��`�d�?J�9�'5���`�'���;aR���9f�����?��🼇���t1�glD#{G����4dK֥�L}���4�&}f�ks�	�{E����
�N���?�~��˖٩�����wN� a��T��XE���08rT��Q��{Vz�
�/U�<�#+*a���U�/H�����K���.��"���� �VJ�d�/otm���U,�w� ���lP:�o�� ,��]�+�/DW�Q�����tHFP_TR�"�6V�sHj�t�m-�(1g:�EI #g�5�bg� �.S��GG9�Or� ���"5�]=�N>�Ao������9�3c��D�uh����)PaI
;�JY!��D�AL�^t��x��T;zb*�Ūz�W�N��P�~<��8o������D���\].y�te�{6�^v7C9AV�̺���f�ׅ!/�H4-�j�nٽ%�:C��bh £j՘��M�t,�\���$�A����Ճ���������S�0�KZ)�K,~.��H:���w!v�U3Wz<�0����G2������ݺQ�U|�$��d~�D7t�f�D	R/�R�&�y$`r'�[���t�
�l	FGn);�1���PJƊ�~qޠ�9���#�X�\�_�#��܄_�S���8�jO�^K�e�5��}xMu�8����o�@�?1���R��	<���<D)����q��#�m%ސM������~U�"��7���}"�J�nD����5)>�zFg�G�ր�7�s�S� ��wiB��ٵ�#ʅԅ��iT�3%�6��Y%�@?��7oq*�&���z@#�f��a 
��{��7- �${}O��uo�[ 5'}�X�S���d�����v���d�L����d,�%��n�ch܏о�([��y*��?��)Q)�(|�e�e����u�$�BfO�;��Bu�%�{�h�������$Ҹ�E�^�aد�B��C���"���H��oۢ�q���\��oqYү����p�ґ'�t���9µ��8p��j���t��z2��ю�$0yt�m鶼*0��ې��.ó�R��bt^E�҅�>M ��Ʊˍ<��	�fz-x���žһ�'����B)E@��9?^����_�*>ES�O�W���2�P����hE�F�%�@$��:�uy_>��Ę���\�B��I����E�&�`g���[|37��UcU]�
[�E�\.��r�8��lsak�WvQ�]XeZzR�"��Ög�����ǵyE��������˗P|`Vq�(�KǙy�5�-��a��+��N����{n9�5�o�X�;_L���	�F!�y� �S׽5ú�ݒ��l3����T� b0r��
��(Ų%	tUh�~��9������{�q2|�Q����HJ�� �P�iz�&n� R� AM������d�wz9mx7���4�Zb,;ܺ�^`­���WNc��P�Q$ܕݟ��H�Ks�0Z���aFJ��HZ���O~f�PLe]��x��HsZ���vu��T�U`� �j}چi�4�4�^-@��y�N�|��?�p���7]�VȈ4.D@�*�]O�P^�_�S��:�m�2^C:+�yO�d�~c�A�D��/�����Z���[P�t�8&�R��u~lqA�ʝ��(bO%ő>J~%aY1���_3Wڒ:��܋�tN@�� ă�H���գ`ŵ��x��T�<�tP�z�����.{_�G=A��񘆙������e��{�����!�4e�������暕Ar��|^���gl��ksr�2���Ԉ�Z�\2���B���%���=�C�
1�\�͗�ѭz�d���2�4���$GF#V���$LY?#@�C����m�IڇfEoM�����U�إ�ڼؘ�p@O��]nkxv��/Mp@v;HJ8|�.U�.0��J��Nbn5��TF
 ��?(��7ǝ��9�?�E>�y�?�-�����	�2����3p��y~u�mXF����#_(:^(�{����yF�k�8"g�Z�:M�G�@`!ȏ�_d�l/���i�9t���P�w�A!ӁL0�󗖎�<�8��򔊧�����U���C���Q'5�]Q�Q�ⷷm�ð`�F��9��t�փ1^?ꍦR[O�Eǋ��L�˼ �s��W�Hgs��Y��>����:���Y���W����Q{� a���o�6,n_)��
�79��襖���~�ۈ�B�gX�@�h��Yy�����>%'/B�;~>b,Z�^Z�U	'%��fp���[|�RȊb�4��ߛ����S/1"�,�[l�MH����\3%�"?|���@'m��#�CT����L�� �mthM9!��(�$ ih��)�T$%A�@ɼ��e���[����6�\�~�b>�K�kɫ^���"�����(	ٿ�'^�)���J��ſ�]��>�^��	��8o��㒝$����ޫ$C ����e��"��?>�;�#�f�w	48�ֶB��������?��|x����� �0�3�a�$��+�.t��/�x�$/I� 5����/�IFp�7�I�\�2�z�j���x�yc���dpo��s���J�zb\���'�)��Ց���d�(�+WQ���=�%�µI�5�q�Lg-zDS'�`��l��v�!�v锤���4�'�>N,��A|n�`���pp@���
��� o��Ft ���(<$��J���r�`��.��.g�,O�D�T��e�L�/6��Zm�}�&^ҁ�������Z+[?Ae\��T�O���GG%A�?tMt��!_��+np���ۗkJ��`X-pB��Lʞi�aE�ֺ�F�����s�^d�+l1r�!�!ɉuo�_1��(���/-�5>PI%yq�pv%��S��bm��ӵ,t�m�o�04��d��!��m���7&<2��a�_)Jx/��-�,�m�X� ���:v� *�H�)��G�ۜ����m�~4cx��^�my��*`�PXY�{�dҺ��mk�����S��V����7�ei@j��<%:g/��"i��VJ��ӌ�2\?s,��k]L`#�$�Ml���4n�}�
b:2���̝,�>�CL���(nl�ԫ4 ��K����8�]���"UT�a��ܝ��"�g�w��{v�@����0��Ǵ�yFRV�ɨ��r��x�X��/g�����P�+PMo\�:&���]�ٖ"�����Z����\m�\/Y�!a.�2�xW���ּ�]�"��5�W��P�q�YG�`4+���kz��U�g�>����yO)�hg���v'hb���'c��9��'��� �I�p� ����4���kk�CӼtR7�B�u�9ۃ\TvĹ��>��@���rR���i�����`�����.����0�����p{0BФr�v=���5���t	Q�oC��-{0n7.5�rg�{3ۧ=p&�8�r�l��Ĝ�������ہ�H@��u��%HҬt��{�����B�������oXZ��93)�tb3ؗ�e/T>X�R�����(j�m���!=��vӾ�@��x̇D��59���Z��6��@��iE]3v���L�