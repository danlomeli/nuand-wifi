��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� rā�SZ )����C.��&0C]�-��[�3�-���+��պݣ�k�J�vo`�A�����f����u�X���v�=�а���]Q�Wۿ�߸�=_Q�X����j>��Zw�K��SvX��ƥ.���#�����Z�0���#7{��\S$��@1I�QX~TQ�E��db����۰� ���>0�%�9�j汈��}��1� ��2���h�G��SeY�a���	'<x�p��k�H`�H�j^y�0�s�78+���ֳ�`�R3dW��_��{p[�?$�s0��#�zS�_��bH
�c�p�IL7]� |����Q�� ��Rr���=��E즕2%�����`�^��l�q-�]�p��jf��Ӽ-f%H���ȳ�>��+���M�71��4_�) 3�46h�rb�J�W� k�h~K0�>P$�_n)���5�r�j��W�J&޴o��$>��6��ŀ�;A~<6P��K�~��f��*I
�Z��}`q���ApC��n���g���3��-�іrO�mF���,�$��@�BI�q�}��Ȥ֐����î�䂧��@������U���vU������ �T#K@f�㯁����|95<@���+�-�)�����K���FI�k���*@�m&���
���ma1[�2�u�I�\�U�yu���o�|��2����;�W�W�}P�K>%5�'�8���׫=����k��,�t�M�0�8]q3���N���GvZ�#z�HM���f5�����;�q��Pj����H�L�}��T7���z@�o	%�PFmy�lc�
)�8yIf�o���Z�"4��r���o�6˦��)��"�~���6��}�pY���]��
��K,�	���1D�̹�@��$���(_kk<| &���x,�u��Sm��Fģ	U��U9�k-��c�KU ��1$k�):h�����!�Έ>�l�B2A�V쉀�#� o�Aڐu�Q�%`��ܸ��cb.�����E��&�Ѯbz-V*�E���bnjۜb>W���z�<\UlA"���i��J��Xj݊���	p��k��1O:�$w%�C�\��H��U���Z�W��k�B�E��d��/���|�0�=o�g����/Z^����X@�N �Y*E�M��j��Ʒ�G��V��$��Qhw-J���,�B�����>�n�N9+���̍�)ТP��yw�~2�]�4�E�,��$&�_�������%�#P� M����PA��[�Z]�ϒ=!�ܠ��T�X�`2s��gq�D���&��%�?�Gy���4E��[4�͹��*�r�S�Q�����!P<�g����j�m2W|���i�:�?���_7��[�@k��v��I�������,��u�T�䷏Cë(��5<-�����8J���R�[{{l�Ijt�d�	0�:�K���}�� ��@W���D���&�b�kݿQ<
�d�dl�\aJ�n��En�V���pT���u!=��$�Z�
���Ѭ�!���w�*� ���NثE�_ *X��F�A
^�7��u ��*r�ܜK	���7�,+�iպ��z��<�7��x�j�ԡ��ܿ�bx2w-�lvDd�T���$:�k��l��Mr �n诗�Tcpb������/��h&�=��|�B"����Yb�=���t-�B��[K߹�zKVX�ʳ���_N��hF�Z�3 �<�~[0��s�ـ�`��=�e�A��l1N���������qh��՘����U�*ן^��^}��Ju'ք����[�l��G���p�clB�A�8�6c�=�lꋛ�I�h�8��M����z�6 vB��Eu�b�9�uY��*�Z��v�A��Xxx2}aP��ju�9�t��: �qB��W=7�V�Rp�`����]̹���"0�H����D�!H#Rr�6
�TG0��fC�p]�v^�ѐ�p��%~�h��	��s���o�
"��63����u��*S���ņX	4b��û*3#���6ȇdÄ��ß��Lm!62f�q��yBS��Խ$��
�ҚY��I�xI���F�a�jv2?�g9Yia5{7��go�a"�gF�ư� H���Q���W��Oø(��E�бm�LH��6�M�g�&,����>�3#�sD h��~*�l"ƹ�=��)2�8c����[|��0t�"Y�8�O��S�I��E+	����=�_�S`�GOT���AO�c�:Qk̠x~�zS>C��8����*f�AK�����n�,��(p�QL�5�ٶ_��7�zft��Nˈ�Y��5�@���r�	�D����eިh�RO��EJ�x'�5
 ܡ����5�I_h�� MJ��>$��:3:Q�Mw���*<x�
�v@��fv��1�N� ��<�H�i�L!�����R�ڈH�с�Ȁu�t��穧�Z  O~�mB�=V�`?=Lp��Κ[ 2+�Ł�JG����	�D�/VX蚌��sQ���	y�愼"i7h`�kzٟ�b��]����
4���<RL/�McܬX��u�������:~�x�9��j�#�����4q&e7�R�U*f�	d�W'���P�0�y�)��M��g:F#��j7 �Y�#���a�V��9C�G�+��n�yvT(����� �XCU�?�	��u�u����vق�@2�z�M[��n�YR��w�/�P�Dt��MDι�I���m��*��4���Cs�W���g�.���jk�v���8���m��Ìٚ�{�ށ�,�I{eAg8�Ĩ.�h7$�0<>?੢J�5����5Ҁ���?òs�6#�<v��v�׃�<�dj}�\���%ń�� R�q!I^�#=�~W��� ���f�5�3���Dc���#}� :�H�B|!��)���m��a�-x8�}O�b�V#l������Ob��f�^J7�3��O�'!��qb|X����]�H��5�B��`|U�_N���������� �[#gÆ�]�[�U'��A�����F�Ѷ�;p�
�*i�z��i)f��E9X��W���]������j��60o���������l�I�+�p�ԉ������܆��Y|���qr������Ǖ��=�-Rv
8-�/�rC�P������O��I�a�}��J5�6-o��-���%�hPB�I��VO����ռ�:`�2h�O�ꩵ2|dn�DO&VjH<ymS� L�(��9�Ɠ��2���o��|�X��X��{��Qa�*qI�a�\�M^O�p���m�h�}� �
�
�	�M2d_�w��2Bj�4�i�el�G�3Fl��,�j���!�����Z���~�r2�߫�"J��Hy�!���|k-�U#�P��<f�A�mzpv+�����xr
�B�~��
�/�)L�yE���V�5��EZ���0x^S�f؀hQ
X�R��uq��
�RЪ|�j�,�O�o��"�4�5������+qo��s���\A�'<E����u���*� }X�o�	�P$�X��J���/�`*����KB�CS�i��y�D�38ރ�S��+9��m���O��v"K�w1�xJ��d1P��&��NtK
�׳�P+}#��ٔ��3�,���	��Dk*����*vϾK���m��7f�bLa?�iS�
T�P|�¥ˉ�� ���7�D0�F�3O��u�+���jҞU0k�&yW�瑝�����(>�A�g��(Ugs��}��_�XY�������nA�2��xKٓ\'8;h�0f�Ϭ�J���t����9�����	��`!E�5ڋ�L��q�o�A��e�&W�q)��-����fM�n.�$��������J؇դ�,8*�i�ޮ�1��,��>�Uou�uX��?�Z]�uO��,T^6�?2�b��ϔeh ������	jN�r��J���3P�T3��A��"h�C�����(�^���w�L�D�������$�1ėJ��X��Tw4	��f������CFX{q7�B���#
F����=߈}��%��J�`�x`��+B']�؛�"�î�s�b�n�'хI8�w�Zg�t��1�t����"��wQ���ܦy�P�ֿ��\/˖�����=$?%�4TI�ǘ��^�j&P���w�U���Cg��!���f�<"���:n�s����������d,hv~�RN��D���A2�޶�u]���v-3erG�]v�H'O)�07#t�Vj�T��9˶'i!Q�0�)	q�ҋ6���yc�-����K��c��1��M��'��93�KHR��V47���k	��zs9'����JSD1D/6r�\&q>N����W�)+Y�W����^�k� EuY9�>�p��� �w�"r9��f8�!A�m"��u|��)��&���ȴ�L��I㺼�O����*��u�͈���ҸZ1����j|f7ےF�A�ޣ}뻮�ɡ�:�{�(�'}�K���̏�Z����)vt���]TB.;a�Mق��	`���HWJt��)�SvTRn؜�0�ㅜ��|X�qu�&J,�����ߑ͐&�8�7�o9r�'�?ևd���;�0&5��M�Y�r�[����u.ۘT����6@|����&������kT��f� <�DN����g�=I>�	��6@l#" �t���D84Pl�lPwC����s@�h�U�M���\tb��J�u�1'UF��tg<j%��q�b�%���5���*5o�$G3�¿}+����#9V��C��7�4��G�,��z4 ��e�\�����7bWdO����zD#����ڲ�;a�%Q,1�sz�!l�ѧ�yX���|$t���o1�����/��3o������h�KRY�!0o�m�uv�SG��ltv��r�hM�'bҡ�$4}�|����K�+�-��QsO�Z�V0(�@]L���.�n#��9��d���e3n�RKt⨜"<�~��!+KK��^��q�����S�W2�/�6�$�|̶Y\8�
b�-Ev�����_�~�k�.�=��S��:<�ܬ�c'q���=h^j�2zE�$���y����"9�-Y��Pief���ga���.��w��D���]n��A;s��χI�[92��!�)"d�<6!^�d1EZ�l~C��=�n�BR��9��8%4��=��'���{�9�\�)<y2%
/|\M��Gp�'=u�&5��&�11Rb�ij�6��X-���A���z���;q���'���׽��^p��������]�!xmy7e�(�+#�Cc����ng�QН�y�T	�(���C�a���!��r�e�#M��ط�|*�ZA}>��� �-!'`����'u.�x�#��*��N�p>4��f>��-H��5�41���<��l������m5�V��/B;��$�G��vN�Ҋ��$���d�>����
�bTY��M��M�:zH�j���'[4^�Z֝��.�����$�06��\�|o������ ��RJS�r��?Eo�@l��b�:]�X�4�:Ft��톌Gg�:��ǂ�)Ǒ���U���=/���%�)�8b�����ނ�-yqW��D�c�� ��#����o�/�n6V�.~���㋳�N��7�_!]���;�73F��dz�I�Z���FLE���`�1�dX���:��;�M��8�KU�r�]* "A�'T���oT'}��a�� N;�k���� ��'��e`���2��{|������Ԫ�����#�h�°�"m�"���Hk�m���z� �5Os'#S��`��~�w痝���ޘ�4�h������*�7��F5�%E���%����	dp�Y�kse\Ϻ�=X�[�c�������f5���7�J�hH��`�Q9P{�l&���]͠��W];~�r(�֢�{��͔�������,�2�r�`���
��B���rVnw
�UB����ٳb��@����Hu�{����a�Or����]"�J~O[O�Ay� vބ�`���r��]O4���]Y�K����i��k˝N`֤w`6i�*��~U�j�(��~̩��қ���ݽ �h��fyK7��ͱrrNk3�8:UH)�KXp\� ������S����I�����I��y�F�x��^�����=�|�u�_ų`z[M�o�(f&�����0��Qo�lo�)���}�F�1Z'��]�u�#�x*:n�����M
ݓ��^����١$�]����/!�4l"���񺺄��ݴ�${�R�>������ASg�������6����@t�v��P����UQ��`R6��qX���ز�7�XjW�B|�T�`���^�]�6@C���o�l�?�D���vu���7:����l�<&��^i����ͫ;��yD�.71_�[�vЙk����R�|:��f�65)K���� _��Bd��ϲ�f�˛i����11Ǵ�\�Sx�
s����w�ă��7Je��)_Ў�j�aX<�扐�@���|�O7�0?xhR"2��r<��'�l�\��]>� �V�p��(2�5�ʕ���p3�h��P�)%�&2L����aLEJr�؀T��uH=��=&`�&/�X/���dr��*w�1�B���2��eȦ�������-�8k�!r����c� dI\g���xa?^�y����3	pE��Z��Ic���ܛ�&�]6f��Q�i��A�Jyk
�����g�^���x�C�#���z�Շ�����¡_g�\�)g��+wu��$(r�%Z�E5�_P.��9�.nJ��k��f&8�{� �wk��```�����D'?(c�Oj�N�Q5��t��f��^������Z��v�كv���:�Q"\���@%��v3|H�J��`�3�75=R�w��M�,�,pH��'Ca'�\O�c#4gEN�GN���4I�)k6���~�^����X��x�2hB{Y蠌�Ȧ�`5�RA{��`�	q��6rl��`�KD��o�N�|hJ��T/w�|�;� F�s�A���_iup�|�:���ˎ䪕8?W�Q�Z��-��T�8m��z�Lׁ���x�r���5�u:s*�2�a�7UM��z� �*H��-�ǜ<:�V)8oC��T=��g����a�_L�����p䈗��#Z��j�C�����`Ce��}�*���&���T߮2:E4��y�b5��a>`�8�,�hE�П�j�,�[1s�{e�Q��@��sG���?Fi�AL���GQse7+&\ۚG����0L@�`:4ՈJ�Xہ��Teh"a.�L�C��X@�42�@
���u��S�[����o�=���%.�0��X*�?>H�`
&Lz��>��M�����`f(߉7NZ����'�.Z/�lDPX�O�����`~����#hU=�]����qBF:��a�\���JG��kx��6\K���3]�Bp{�$��h����CN|?�����̌�2.�_�K�y;/�>�@�[��g4:΂��v����fDT�ܼR�:����g�@w���I$��ga,@��K�u�C+�F��r������f݊Ѻ�����{��v|������G|Nn9R]Υ?��;j����C��^��>4���V¤��m���kT͋/Y�U���q�n{�Q��/K��������A�K�CB��p�M*l���v�4FWp� �.�E�8u�m�笱'=Rm�Ni,o�H��!�����pu��%.�@�ە0��Joc9=�N2���x�H�#��������y���d�4ί&��.�8�BR�&;��R>���@QY�\��}O��P]��5j'������j�a0~\��-����TE�;�2~�	�^��hή����Fs�����W�:n� �l��i�����X��ӭP�6 ౧�Z`��߂���
M�%Y,�E�c2��ߚۉ��/���Sw��n�"����kB� #q,XٹE�cYg�LTR�����`_lf.��.aQ-X��%O���M�Y�W�w+��f�Ka��\0Z2eE�tU�p������K�@52����3i*]���|���[�QtM����채����m@���T�����Q.����F�XBe�2�4vq����+�vCaJ�3\�^YF�n��
��,�jy��YΓ�0�L��� ����-���������͟UE�#J����e R���H��}v���=�Ή��:+Y���z)���2�����1�j_vY(+�dO���;�`�@8�r�[��j�m�a&x� �}��՛������ײ{oc�w�_4@0��*ґ�5�ÞҾ.�6]�:��SР'�#��]����f�?�S��Zt�~�FƇM���އ�{B�X��嚊gUU�z��+@��_`�e�a���g��������P.��qN �@� h��c䷬���28��G y���J���ss�P�D�<�sٽ�Km{,rzPޣ�مEБ�8�׆�������!���D4��f��y�U�3��\'h�,X���������D��� 0���R/i¢wd}�r�K���K����<��KNͪ\9��^?5HFU��ԫ�\4��^}%�\�|Tm��1	?��q\/��E�@9�l؏��dK��1Z!�8����z�R�i�A>�s�R(���T��"m��#0�@]4�9��Y��l�6^m<h���f1ݍJ���l,��.+cA���Lw������e$b���uJ!	�hO��ذ����̯2��������� ����JS[r�o�*L���7%����1��R������z"�E��ן�G��������H�5W�vÂ�n�&݊����J��2�I�Nժ<���<A��o�.U�
�TI�O(�؇8B!*��s�d�q��ˆ� �(�
�#/��£)�:�X�c/^[��@��)Pj��wV�}�����.����@�e���]`��Sȷߕ�1���6dQ��RŐ��8�Cuۄ�:����I��Aqpݨ��~!�M���q�}��e���nǘ��$Ǝ����؎�80�H��� ����_o��}�@�t�0C�I�H��3
1I�c�␏�ݱ
�a{Xbٸ�g���U��NOz�V�(�vC�m����ڲx@*���=�c][u���S�sN�?�Ps���w`Pvh���R���8���	�-`󠈩�	�4������V=���ΰ�U�M�Yp�(t��� �����b�I�^�D�Rlբico:�	Ѵ�����C����m�'Ne�:��W��H t�C��_.("���l�Ll�Slf�@Kg�{I֕n��mi-#J�I��U�ő�UʴE����(9�� 7��{�ƛ���B;�:#9RY�����hU�Y�2�?���Ǉ�M<1{R-�fT/+� �e���6~"2��x*!���tU��c3G:��Wgmq.��k�q�A�f�X��{�������f6
B���j��$�A�1�R
���%l9�x�h��9	��� �Ji����'5�:�a�� TW�S��ҵ�>
@pt47����zR��GMS�_�@���6j�2�'�U#�F�!��Z/�b��#IcҀ�F��rI�Iԥ���}�3��/7x ���:2epk�:��pj\�\�K��G��	G#{�L�t=j�%���߁����B�Ǟg�J�t�_�+o+ć���6KHA�1����Z��gSp�5P�h����K^���$�׬��A�&���e��zi�`�)�"z �"�z�0�6�F��r�Nc�ką:�ؔ`|��d\�1Me��@z^3�Ig<�f*��F�������������Z�XJ	 e��������[�/�F~�˷�f5�S��y0ٛP�O8����iRՁ|v�P|�4S�鼁��*o!m�q�|��CN�4��{�Eq�ad���&IUP;��sސn�^4)��mx!I^N�)_�?YK���UZ�#y'���jr��0W-)�G4h�+�����7x��V}I~�B��SB���n|ʶ�0�R�=M3��W;#�U�)��]LJ��>�aN�����lIG�}��q6]�T��>"��gR��N�2�[M~�9�.��y@��.�دʂ,3��n��Y�Jh��K��L���R���𝲺*��?xi��EȈx��*����.�J@�_��o�<�f�8z��9;V}�C�NS�e�w�O��v��Tx8��ceߢd&_ƅ�~��z�f�k�?�H��i�:��-QϬ�v�JVG����e�P y��yFr�
�~���^9C[�A����b�Z71���W1��R���O�+�g#�wk�n��t&�h���;����U,O�4m�ps��9��	E��vo�z�4_�}���6dG�x�4ɔC0��-��*�ܧ
�eM�N���lz���/`;�]�Џ���<�<8��`}#��Lls;p:l�]O�u��ső_ +/wB�2�g�μ�#���/w��N�kX=�Ĳ�sueCu|���z��:N��F_sI"�\�L��d}��&>=�Y��"��z[��}�I���j�L�ctd6�h���Ɓ���PZ�H�a�k���ƨ�̥�f��*�ǃ���#�sOr[�a�K�R�������1(�R�<��$��z���K�2�C����9֯{!F�C�������Mw�� FKD�Wv�G��R-�V맭8~Ǖ�[��H�������� �G��X�J��_3�#1��ɳ�ɼZ)��N�tL���f��X�.Z|�ձ���YJ��߅�kw|M)Z�p!��9=�G�^e@Ҝ ��GꎼfiX�F�Rp�(���F@{��l�ڄ2�b��yꀇ[6��_r��F�p(��n ����YP����t#Ȍ��O�i�f@�nD�U����_�""|V��:�O�*�M%lX�����$��v�T��HL����#E��Dϧi\ԛKl0�E5�@^
<�C�%�����r�yw�$�������=����跕L3=��;$���}���W���M���`�����0R�1���{�2rue��y��n/�͸t�B��`��-��y�o�ռ��R�wt��H�Ny�N߰��Y�.f�d���a�����aY�)��2��A+�Q���iF˜Gs^s�-Js� �Sm��.\L�!e��k��2
�I,!���"��ޞ�B> �m����	�����Ҕ!�j�n����UN�by��\X4�s� x�py�!��u����3�&
�G��-uU�uG�0�L�II���p��UO%ck�*�������/J���.U�O�IE���h�s;�|�$��!�[�>���|�I�R�-��|��ͽfɠ�2�d�p�E�,RT^�~�C�_y�$�7΂�>� B������ɧ�J#TH��4u9����p&n�������ixw����:Q���&�\K��\�w�k���YFz�):-�(�!	[��*�,�ź�������\���AY��о��v ǵ�5[��xQ�l.����u�r|<��N���NH5#�s3l�0�n7|ٕRH&H@x��nGZ[�>cԱX� ǘjE����漢���1b���OQ�g	�t��9u�n���u�^��	��I+޶�#HG�9*�.*�xV�.���׏��:戥!�0��#P�~1�dz�>�����~�a���i�����w'�(��&��9����i�`�0愼�g��<c�`��'���;�5ԧ+��5aN/�97��PJ.pD�T
����zt'��i�P���ÝDD�iذ��f���u?�PM���~�
3e�VNu!֙0]+S�8�Ѡ<HJ�t��־����'
��U]����g)�W�s��׆N��|�������.ວ�wX#�,q!���!��g�$u/M᎜�S��O�}�o�T��to��bt��h �����sS|��4�ܝ��ÿr��&j�p%42�րkXh������j<m��B��*�ԉ O��%��} �5s��E��>�t?gߔ0U�JL7�ӎ)�B@g;���e���y9J�J_m��g+�:t�~�܆XI��k�y��!�����b$��}�m��IVA���mE�0aN���_:3ə���M:֥��M����
�t*���^�����$t;Y�Ԭ��D��d�5������݇u�n%��N��3N�'Diƪ�)�K�H�W��B�ܥ�G�����6Nܙ~zϹ�:�R�T��R���x�:AsFR�cl@�����b"^>�6O�z�Ȉ1��4���~6�q�I���
���-�x�g���J�cL�%���9B#ز4q `歳��`ۡ�2���x4ח�Ԩ�"bb�������$�)uy-����+�B#�Y yx�߿�nk��2[,{8�>y��֕9�����FNq�����T(��<5@�/ZEk65�ҕ8�_�Qf�%}I#�Me:ͳ(&#V
hذ+�{�u���.��{�X���t)��4��񃥷u�)G�����ӿ�l��C�a%�)Ӑ؊�G'v\쎠b_�d��P�s)p9��v2>��W�y*_�n�(�q����
�̹���,�CP�8�z���;���H���b�J��?�ɚ�H���x�Ic,�{q%��1fN:�Q7�9�#��Q�`nv�;���)x.?=�˲�8w9up|�풭��rIMj8�R�V�Ӎ��>3��b�T��n���9�G.��/�si�c�"��=��祆��p�_�.3��a!*��q���ofB|�ۛ_�3��l!o��!,#��l��B�`��\0�2�h�Otu],�A�Ǡd�cB&���oАs��l�YZ�S%-�Y�a0�^�2hH�mO��I>��p���~�HQ��d��RU=i?�)���
jg���Ły�Ǻ{%G�z���6-ސ��E$��7űY��3wz�)��'[��Y���^A�wJR�b:4Fkڹ�!S�|�U��S
�^��y��	��aF����S֔Rj�B��u(VI��}��'Y��h��P�J������R�kDrh��xnMJ��<�춒,�e-}gٿ���G�QW4����3�Z,��PJ?�'�����a��ؾ&�%n�2bn����:)#����d�ce���y�����0S�Tfv���	˃F�������~k����ͫ��l��Ϧq�6����.Qrem�P�,���$��A�=��P���vj��2b������ԁ��n�-K�o69��EG�(��m�	!�ћl��>΂�i)�ߍWބ�ڻ���K)�ÏQ_�s��7_td�"���/�lLC�˰#n���E�_�PKI�n5!�\���of�8��0�%� ����aHg+w�P圲����� �)�l)���tw�3�Mm�ی�g�j�:��a�	�Uh�����C�V�_�=�#�l"fD�Msù���[@L�3�,����O�ظ+I��>�R+T�b��9����-���.h��2�����Gi��؋nQ� ґB^-�R닢R`RR�Cv�?W�+8ȹh1ڗ����c/ VH���[���ىMv���1l�~�Cf�� V0����rS!-Fq��I���y�!*����#�^��O��=��Ӷ/�=�~���- �D<�bb(S�V���-W�k�{gx�Y��ю֔Re蟲����k�1�b�N�!8a$��:�Ъ}!},�+�R�+�	l�@vHj����[Ǆ�P׀@6��<������yِ�2ga�gg���}o���ڇ���S����S�1J�<̞�Z�n�U芊�)E�r��6]ڋ2����#Z�J�uMo)�!6b�7~�%�&d���т)��}B��(��5�"�ذM�#�Q��
����*	�����JLH�F��N������6�qŬ���E���e�y9O���,�4��"�)����A%�ʵY�e��#�x�C�_���ki����|�`Y�Ϣ�7"�\���_�䥨����#���F�W�����C<U((�Քor�i�4x:�����؃��
Lᗄ<sIrj�C�/Y5Ӆ��jeR�+��!�;p������Q��K���X���hHi޸W��Hvu׎�C�R�������#�iqZ±t��+V�J+��j��`�a��(���ϖ�@��cX�Â>��E��:��A�����}��w@f�2hkz!���F{.βb>��u:F��&`EP@�  q�U=ŻkT�0�BX�%���&���yf�:�dOD������@���c$�-�=��=U\:(H��Z�4�U����gm�1B�cT�Y�o e$�8��}3crY���b���՞���{�K��
��ݟ� ��B�7�7qu���Z�-��<�;�<\.���>�����A7�+'�,�k~>S�?�f.5K\��R�b�Q�o�p�'���������_4l?t��Sd�[@���	)r./[zi���^
����>F\�	�f�����e�$�5i�s����暶3"{�N}P���6͢$?J����Rz�1Q¢�b���$��B:jׁпCȩ��l���Q}�s؆��j6�`��^G�M���H%��ݑ�)�+�o�aj�k'MK��v��̯�Z���:y��b�ɶD��'BWs=LВ�gm`ɞ��;K�̥-�"G1�Adm�دZ���6V<�1TP7��~���=��R��mA9�n�t��L��_x��ʀ�����vx0��X�$�s�PD_�2�vw^���G3)�z-�����}.�����Y����;�m��0,@�ҹ!ž1@Y�����O�6����蕈u騝�QC7z+��(`ӣ���W©��ɑ�׭'b�C`a���}��<��VpI=Ip޺�`.�*��U�:�����m'��>��- ��a�<��Y1�7�g�,҆��s����w�}�/��������t����T��G�^w��څTf��.I��*����a������Ӝ�Dǫ`�j�b	��<F6��\�p�jc�[����8�Ŕ^'��iZs(\� 8A�՝��&�$J�V���$D��
j{�E�%^ѣ@��P��q�n�Ҟ�c���r3�/v�	�/er��2��ńF�G�2³i��L�	�ȁ�
�q��5��x�O.���)yn>����샅m�g��ۡ���=Z��o~e�=�a��Ji�J�s1	�_���V��4�C=���6Z�7�7K;SX,��:Ixd�
�Fn�ђ9�9�a�k2���_~ѹ�3�)<�Q��ߑ%n�6{v��JA ��L�l���Ya����EQ.;8/kk��S|��&�*:���y��M�oؙ�8	 ��VaCi�w�9k��T�ނ�C�gM�YI���ٞI V�N (˖9��#�<�����mr�N�1/��F+&�ڌ� ?�Y{�(�L��}
�"�w%Է�����iD��ww2ܫ���+,<p&*.� �G�q�'cO���I��n���Cv6��J�5�^�H8mk���H>FpDb�`���Dy�R�Wh��up2�u�����Ɨ?K!�0z�ۇ{���F
X�9{�)Quh�1���k��#O;�|a�5��\���t`'{,ոv�Z5@٩z.U�:#�t�J�W����f�>+�eNC�KC��P�u۞�b+����|� )w+��\�G���<�&��� d��O�l" "j���<m�5�Um�=/aI.�H�e�-=�<��fį����_�P���h:�xU�*A�|=$�t˾�#��=!���X�>��F:��~ҭ79�`!X�������A��y:���b�o߆ߖ{"��6�GiL��X���Ԫ����\��˶��{*\-Y������4vh?�1�s���>G@�69 �C:���.PmX�5n���,�(h�=r����͚�cᳲ�r#6�bfIT#_���:��_�~5��ٰ�ֵՈ�%�����ۃ���W�D�xe��gu��qJ؞��E霡4��u2P7��.�&��ql�U�'h'�q��8ArO����1��&��8<v��t�n��<I-�
}�f�}X�P@}�⻆F�*�rӃ���bP��'eV<�ԃ�}gN��eQ��\O|��e,�7jQ�&�y���&�0&��)���>ރ���4�S���6x�eo��8��]co�f�	����U�N��ݴ�Pڭ�䟬���h�
�6��U����	��U��z��M�׬tj	?C�̄R�g�Iv����#�����,�ÉK��x1[����a�6�v�坐#D���	PLX��Xn�́`��Vkub4��W6�?Dv"���T��P?��t8�c��ە�!e�� ��J�TR����g�t+]򹀒:��� ���螉X�X�_�
)牦]��Y���gzT)C�+���)��z�ȏ���y���ͭs���H �l�w��������6�'�ґ��/;[�z��m.ǌ�e������+�����6%�-���k��{���2�䂂AZ�A��i�,&�X�l��h|1>�}%��5s��<@�1L�#�j�'�д^�>�tz�J�W� l�{�h��+����og4�V�\�LU��wI{uݹݓ��gۢ�I�:�-�-�ٛ��v�dX9eK��}��m��~c�`�nL��@}	��N�0�b�����i���{{�zÐ�nuk����#�G.���薞��I�U��e<(���/b�Ll�*>���`�R!6+�2�����@��4������n�daZ%#�[�0��\Y���zd���P�N,�y�;Q�K��q���m/��g�#[���Ϙ�D�������8��͙Э�<�.�T�BEѰ�����|=�ęF�uQ\��	���Ah鶻����"�J��d�f����z�2�zkj~����m������M���g�Y��f�)����s)���0��%^�EK����16aW�$�`(n[g��DB���HC(�{��!�w��Ҭ=��}���}����8�x��W�͉��$�V�s8�v�(��`#�5&�%_��+�N��F6n�˟5��BZ0rl������KDW;��S
�m�X�CB^�\�X�L_����8�������K����$?�tn=�g,.1��WUi/�H��2^�@ :����i^s>X�\��@�X�h�z߈�������#�ʼ4 _��+$��̞\r��/L��$�xM�Pl3B5� q�l���W�TH��ɣnթ�����K&�x����dcm�k~�v�7��Q#������f~3�����~��Ȝ�x�y�.Onˢ��
�go�6�sK�pN�W���)u	 0�-I��!�xQ��:�{j ��w�	@�9{���dy5������+��~�ȍ&�SPTY����0��Ep�o���k-\%4��)�/=��˸�7�\ۮ�Uz�J�ޟ�O1^|��ɔ�~��\	��Y�Y��	�m���Ա��
h#Jr)���]�w��q��5��z�F���"t�q�V[��h��!ܹ�Vk�;N����^���o�ִz�؝9Ȫ���ja��Q���w��;~�&^N�,Mt�8C�WTA7�_�'9na�"��_�~�#���
Jz�4�;m4)�D^�[\T�X0��NM#1�'���6�0��2I�ś��^��wC�(@5Y�Fhz�e�Eh�aY�����er]��NNN�xk�X�b�������D~U0mSc�+�;S��0,O}k��S$	���_Ji[B�z�Y��c�{�Оy,٣=�^�I"9�m��L���}����ݫ�3s3��Dw6��3(�3O�֮'c=��3̴: O#�܈�,�$���r��J��Y�P�|u,ڃ �%�IG�5�?R����_��H�6�'O�h�׺�Z3|�ʊ/"�]:�歱ή�%nu>�o}rY� w��Zh����h|��-�Z��j,ߺr�]p�x��d8rD�\C/�9���_��[�5�ZPѺ!�'�{�{�n�_p�+�w�m2�Gj)�&mc�>����V����YlXܽ�1�5F!�7hg�&�Ir.�3�h4��L�i��<~�_��,�'�=Ln�E�u87���5�r��y�ߊ����X�; }V�N&�FJdW����Cޙ] Ej?rK��ެHgc��˛�#[�j��_d��d�������	�:D����QwEv����y�񀦵W�7�0�f�O��xZ<��D���ee8�1z n�[M�Jci�����h���`������b)�p�+�$E�>�c3W%iY���v:p�V��+N�4a]�)$�kV�Ą�@.�yht-]K+���[N(jc|O�@	g��>���{�i<z�17��]����D돈���-ju@�y���6oa�x����f��=
��=�qY�u:MvY|�v:\K��<���-��"g��_b4R�XH0�h�F����=Vڗ�l�jR,�k���5�R�W}���RM�������쉗����l9{Qw�x�\��ߗ�釪aQ�Hj�'�d]짢3�ԏ��H�	���t_�ָ�B}�m!I�@3�~�ᗷ�{�͒��Az�i
���#?r�%�7���� �ӂ�$-����|I{u��!�k�O�sr� �}������\������$���#���^F�L�jw�З6@�T�&:�F�PT'R�mZ�uSw��)|œf�����I���a�y��,�O���<W2O{ӂ5W�pE����1���$��OQ MT�w�*�d�O5'ws���T�K�HI}��b.�8.f��gY�ʶ���M��Ir�� �D�K�w'���{�o�Ɲ 3�P�qD�k�6�	QO] ��e��5�E��e�ܓ#�-��߰����[�GP��0G'VE�/.�"O�خ43jUnD8x�Rh�MO���5��ߡ�8��b��]�Pl���r�x
�?OrZ�M��p�[��j��{��*�O_�'K�&O�A$<_D��N%�g��}�ͳ.�JO*�M�ēx�uI��q|.��P��Л'b:��D�a-�ꉚ�;淰U�>��~R����R=�^��� 8���3;:(��lA�|>��j����٠�����g��#i2�L��3ȳ 
��*>2'��=kA�m��Θd%�l�ZL����j1�`%��Q�W�+F��@���'���B]RDr�+�C��:&�ߌ�ڜEV�c��uq��w�6�e�e�Ro#x��������=o$���H���F��/�n)�B��2�WE]�2�~�=K�2 }P��O�m�P���^�rJ*�����2��l��tdZ4<��.�9r�����ˠ&�7�|�h�������\_\�Ux�g�".�P��z�����R�ߣÑW�s��Cv.�'r'=1�����m��:��kＴ�I�_��cn�r����[��~u�Du�O�S�5��-������6�<�0L�l��ǩ�e�cSk�������R�$�=ٶ^���3x8�3�Hў3q�w*at"wM�Ԣ�s�:�{����,m�L�x���ۇ4�Z���[Iȗ�vj8^F p�f�R/�?+����w8�.y����]��d������1))�p��1kzZH5�Ī�Q�6���M�l;-�-C���mFnȿ��% s!o��?��?6Z�v�?��E����ʦD��ְs��Z�g��񃑌�j�EW�\k�a0�K��U򩣝w���仗��J�n��pRNo��Um��X�v ����?���2-��V�:%���'B_��@$��ȫ�P`�-���z���S�p�
>����6`\SU���=]�Mx
��B��Me�&�g���j�(�9\��w��3�1A�=!?bm����f����dk�3���Jo�z\���^\~j��]`A���D�OHB��O��	��B�����sf�!ђ	���~*��SEn�
�g�$*�
��2�����zl��*��[�J|���_h�(^�}�^�{N5�>O��*�lo<��<�phgWg\�g����g���Je��1��b�2���S7ɕ^N��f�O��w�\5���y^��܋�p^y����݉�Ą�J�d���g	�@/��	T��\t�bb��7�/�Q56����_��\fuZ:���E���5Ln�` �s�T���	��;���<�ynj
]=4��2;���9���3�L2���y�O�NhxO��KFSK1�է=��w��tH>t�J���G ��z�OdKp&�6/L��� ��%����@Q�6]Jz�^|�'r��e�m
�W>��Z̓2w�v���W�g����!>��nI����o��Q��L�ϸ�S�g^��C���k� �@�2S�~����)lָ�Rd��_�[�'�ԕ(�a���0D���y� ��+1rC�^��9�Q�~H�n��Z���5�+9G��F~�����sM<�ʠ���`ks��"�h!Ԣ0"�A���}��	ܛ]>q0�Z#�Z �����lY��7!;ٵ��q)mw�5U��qK�A�P�U�B����T���H:&��E��6=n�JI^��=&nB�c�Oy�-QΎH:�����p|�Z��!Izm�?�S�[��q��5��8J:�V4�21+�?a��J�)	�5�BE��Z����gX}'4ݬeJ���+w��L�Jǉ�Y;���	����j�&\����27#�M�m,�EQ��3��X{7y	�b��_W�*�oa�2�l��;�p�:��g�I�҈t�ܐk`5:[_'`!{��|Uy�R|�Y��=|��|LzZ�Q�蔱��E��_g5���`i�7��(���/*׃̒�A���V3}D��[��*vi6�!�pe�\��	n���ȯ9}Z��;�8�6;R�'+F8k=�P'�X�J2#�:�l���� R$�ˣ��; K.KRl�z��UN�FE�e���(V��,R ��A@�@���'(��/����Sݽb*`��#j���i�O/��`ae��_\����Q��������\�3z��듟����������X2�qŨ~�6}3�LFۚQ�L�	~�Jh{'�U�D�=�����r9o��_A��|#sc�R�O5�G.���j�̗\���G����G���,<�8���j��>6�^�\{a�ƪY��GE�(.��EYR�ſc����}�5���mm�z����������i/�V"���!OÆ��=�gд�?c I��lș��*q�������N��z�~�Q�Y~iY1}f\�QQ��ﾩ�~Kx��x�ns��XEQ4��nh�ǕU@�ت(g1zn:���2f�,�+gӭ��X�鸇�D�h�Y2f��L�
Z8���B����b��ri�=���[{�\�ȠO����I&W�#�k5�b��=Iq��m�4}�;BF���+1t��I��M����M:��ޚ���δ%!���=A^Y�.}:��S��O"��KM���vp��D�Dx�T�"���%�<Yۥ�����d��]۶r>�����g@�չ�8G@��Ibx�2��nzXw�6t%��"1��cDS�3cw�}_8�x�e�����3IK�͗��DU��~�#��_)0��=V�{y o�Ȑ�N��QBR���5��:��q�\�Tu�*Cy�9��j"��G9?K�p�:?ǓѬ��3�[vͥhM^h���KEǨu� �KcJ��^\��T�)���[z�� i� �.69����9Q�V��	o�'.r��]��L�@#���N�����9�JUo-$���k=��?]� v�v�`���s�E�����b�ќN*e�����l��a$|�����-�����V��jI)O:֍"�J+[j�u[���l��ײQ���� {*ې��,;�7�~%Z���T�op��(�)A>���2G�G��d�z��|̦���%��/Rѕѻ�N\�Bm��>��ڞo͍37f���޺�8��2���X:U�ԥ�O�Dcq�����q���Fc�����ߕ�Y^��뚇%�C�.4å�9D�#���#�u`�f�l�C���o�S/�h�Սs��,`��+,��|<t]��;_�=�<��)��b�h�4v�A�=I�M��ߟ�U!��P�=Im-{�iW5���/��Nf܄8RR8Ǳ�i�3�q��e�JP���!6��t�CЛ�Ȼ�S!��="�<|M�1�m��<䘕]��;W�NK�7������A�ڛ�~f�=�N��
�P��bf<k�K8�����A�rh��%��0f�T��B�xt��J�	K�g���J�Ap�*�1���������o�~0�@��9���c^U�(��ȝ� �����ۗO[>d�´߁�#D������V�1t� ��z��zn_��YN;�3�ts�@?+�]�5p�x괚��x��Xc��h�4���@A�o���ȎRLf\L��;�-o������n��}��U�{��3[C���*.}���o�'e����3@hm�����m:?z�ט�?4	Ũ����=Y�e�0�������[��p�<�5���͆臗01����aq�"6�`�9��Ѯ&��F���pп�㲒�`ɏd/Ğ��n0�)e���V��r&�զ���t�k��;Z�Į�_fW0s�������?ߒ4놽��rk-�k/�����d<���j4Bc�K��4���
�y�E��5�j��X�U]z��r������.J��u�v4R�&���%7��k_� ���v�ˮ���,�߀�/H�t@sf#�>s���8!�g�L� ����C̦�f1�p���\H�ҙvW�����F-W�q�bLs��8���"��gVuj���vl�o�ǰ|ϿK�@RM�"����G�g5�~��2��C��7v2_��tT�@�T�ڈ��X��"}`�w=���z�С7��r���}>���b��P��a#���?�A�!�l���YL8y�:�؂��Ƅ��Ү���_p�7�x�^��@>2�1+�"��YN���O][	h%���լ�ۡ�?#Ro���tt�ߧ�݁l���8u�쑶{WsA36�3��ys�K|�`���6Y�ݓ���͂
6��OJ*O�_hN�u�^m2�_� �?V�{-�%:b���1�3bq���ZFb+�����K
4�ݓ���`e��I�	Q�Ѐ^�;ƯoO�������}�Ğ.V�@q?��dv��tG.��wFp���Kn�y?'�҉lt^��^�^J��0��=�/N���~����ϝ�L��C����ό�%��v�Q2���R��^=3�Q��j_b͸��ޱ�BȾɛ�#9 �r�~z�~�n˟����e~689՞��o��e�PnI��=��ͪ��M�<���"�(�����q���wI��� �V����H �2�/�	��?�DӅ���S�m�V��4~1�}�|�H߫����^�v��O�A(��sMЇ7	���e���n���x��j(D��Z�1h�b<�KB]�N��)z-o,ͮ}���Pc"���J���z���=L�W�A�`�'����Ʒ��xw����=���\c0�
Y27/b����G��\���8P��if4�S\ڰ	޵�
vA���M?҂@>1b*��<O�O�A�'� M�L�qٳɛ�1�+��x�o�"P�Ϡ��8�3��N���0*�x�|��:`�B����z��kX2�������#�
Fe�gK�H�!?jv��LC	rf�R��-�`�|�