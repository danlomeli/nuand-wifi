��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� rā�SZ )����C.��&0C]�-��[�3�-���+��պݣ�k�J�vo`�A�����f����u�X���v�=�а���]Q�Wۿ�߸�=_Q�X����j>��Zw�K��SvX��ƥ.���#�����Z�0���#7{��\S$��@1I�QX~TQ�E��db����۰� ���>0�%�9�j汈��}��1� ��2���h�G��SeY�a���	'<x�p��k�H`�H�j^y�0�s�78+���ֳ�`�R3dW��_��{p[�?$�s0��#�zS�_��bH
�c�p�IL7]� |����Q�� ��Rr���=��E즕2%�����`�^��l�q-�]�p��jf��Ӽ-f%H���ȳ�>��+���M�71��4_�) 3�46h�rb�J�W� k�h~K0�>P$�_n)���5�r�j��W�J&޴o��$>��6��ŀ�;A~<6P��K�~��f��*I
�Z��}`q���ApC��n���g���3��-�іrO�mF���,�$��@�BI�q�}��Ȥ֐����î�䂧��@������U���vU������ �T#K@f�㯁����|95<@���+�-�)�����K���FI�k���*@�m&���
���ma1[�2�u�I�\�U�yu���o�|��2����;�W�W�}P�K>%5�'�8���׫=����k��,�t�M�0�8]q3���N���GvZ�A����^�Љ+��֍$�],ȹ���{��v���C��(��B��	4^9���Y���e��^�?����麑������<�TG�J�)��кd�1��H�����7�Y�(cd�GO��<#���1p���3��2M��e� c��������U�w w���j-��G���$��f�S�s�;D�O��lӡ�$�i������+抍�vI]6���sm$xt�>K&d2��_j�,��u���G�����&$�,᝾�����5�l��	+�O�7�o4��H�S<�/��*�3cU�?��9�rH6GAu1[��,��Dv	�?ہ�&^)���&er#rL��N�>v��rb�P�M��[�j�a�ǫ������mf�G\� ����h9^a����'@>�]��,�p;:���V^`�쉌F�}�`�z����?>�C�d&���u����ZX���'G_	�֡$'� F�`W�N��|�2k�����!X�y���j�x��Xj�+(�~��Qv����.1I�Z�Ak���Iz�zV)���C|A�A4Z�z�����?�2ݝ̀�9=�h������l>�_��8ۺ~ �벹N%��<���<>*��hs�ߣ�'[�v�W��� ��C )>\����$�0Usn)��j�85 ��1�[��dp�+e��m���������T��4��N7I�i�0�^b�4�g���uQhF똷�E�ޱ�6 O�"?礑Mw����V����l�z��*�U=���S�恳%��ɨ"� oL�=&�m(}>�%��n�ْ���z���M���K�j�`iB����Nʝ?��!t���+�)Pť�������_�|+v�F��q��]%Q0��Ruq�`��L��'��v�I?������J�׹�c����R�I}t=�;n���A���8x�#Y����]�l�.#2�9�C</PS�m}+!02>y\�hcc�;���}_��L�S��⎜j{�n�U`���}�K�?
I��EUV{�tdSp&2�xpBlR�Y�������jC*AH��3�BQ�^���bB��2��9�%*�ݪ&��-:)��P�:D"{����F�q�uV��}�v
3�a��@I� �4��/7����I;D�/�E���f#�-J��vQ�B��8�q@a
oV� ��!��hk�[��	\֮:�Kn~e�k���0163�{8a��^��e�fN7{�V�/J$��#����L�*ՠ>w3]�[�d�+ctl���Q)�(�3�GS�Y_�@�h�|��@㇬��#�,¦�����E�5f�;V�{!��_�����|Ҫժhp0�����ž C��_u�O}uj}���M����۟�tU��Z�a�2������;E��V�~<���%b�9��M-��֕t�3�[��+�Ձ6lw��ss:�&f��)K;�Y�� n�E�b u. �&3�Q��Cs������+Qg�a��e*'&w�6+#0�c��L�ʿȰfi�Di?]�������)���E�9ߙ_�j2���������+���>i."�#f�ŷ�>[��3]S$U�y��(ݪ��S���"�F�w���d�
�J#�?_�[�l�aV���C����arL��`j�4��?�n/�oa$�y��G��4�X�W���Q����L�n��j�SIњ������@/��)����ܯ�!C��y�����/_+������|�H����E����7@eA�Z����g���	5���g��or&���������I����s+n�� ^*��Z�j����'S�͋k<�l,�.�Sd�U�#�!��$�J*oO���G�A�#�vy꼚ܕ�	�<�$�Y2X��:�$�*�餸@B���@.3��}�����@
��{-�����	�)Ht"��@���;L^���2�|��*eX�@��v���p�iu�IH?4�	�ncJ-V惢�WaOs�@k��[����<{`���Lw�ĥg�L��v�4�>;���3���{�\F�9Zo���0���v#p)�Sm"L3�Ri���}{X�ܝ+��~r���w��8]*>���S�L�~�Dx�A