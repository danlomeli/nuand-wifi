��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� rā�SZ )����C.��&0C]�-��[�3�-���+��պݣ�k�J�vo`�A�����f����u�X���v�=�а���]Q�Wۿ�߸�=_Q�X����j>��Zw�K��SvX��ƥ.���#�����Z�0���#7{��\S$��@1I�QX~TQ�E��db����۰� ���>0�%�9�j汈��}��1� ��2���h�G��SeY�a���	'<x�p��k�H`�H�j^y�0�s�78+���ֳ�`�R3dW��_��{p[�?$�s0��#�zS�_��bH
�c�p�IL7]� |����Q�� ��Rr���=��E즕2%�����`�^��l�q-�]�p��jf��Ӽ-f%H���ȳ�>��+���M�71��4_�) 3�46h�rb�J�W� k�h~K0�>P$�_n)���5�r�j��W�J&޴o��$>��6��ŀ�;A~<6P��K�~��f��*I
�Z��}`q���ApC��n���g���3��-�іrO�mF���,�$��@�BI�q�}��Ȥ֐����î�䂧��@������U���vU������ �T#K@f�㯁����|95<@���+�-�)�����K���FI�k���*@�m&���
���ma1[�2�u�I�\�U�yu���o�|��2����;�W�W�}P�K>%5�'�8���׫=����k��,�t�M�0�8]q3���N���GvZ�i�+ C�e
��Ќ�S�v<%���q��e_��
�k�夞��>ZO7E~��5k�TW Aod��eE���G���ɑ-'���?�G$����ќ����8ɸ+ 5ʗ���l�d��,�J�
�^�3b,�����J����#n�zK����z�&��;|�\�^���'e�W�����">�w*	FO�Δ��v���I�h�*�hF������$�!�^��z�;hd��zޅem�g���Ǖ !	$��s���;�j���}�_�vb|���z�YR�c6������ē�o%����li!�M�����l%�]���]� �}!_ ��ś���Nuh�k�)��JS5����I=k���Wlt��|�*�*6�P��T��L)ǣ�6�>@�����	{��6Q[G�����p����B	�t_[n�$�4q!�\)�0`|�Өf�b��L��C��i���C�ܦ5�����c��{��1ni��(����ͼ����S�Ԧ�c��/mW�6����]3C��y~h��:%VM?qE�l�|�N�J�}�����7gp �O�ߥ��>w�*<�?�	������D�uӅ�_ո_��V�+Ժ�+/Tؼt��X�
4��8�B8����*��PL�2���F���fRm���P!���f�$-N�{O�;��〙Y�ZL��^(�`o�C���D���|�@��a�����ර��z����z����j�I�xq�ՁHd`1X���U���Q�8����y=�15�c�G�J��de5o���U%���Y�uuK#;G�����Y>n"y$��U��.���4&���Z)D�`|�Kd���z�Z����N��8F�ũ��X����k;�����;����y����S���x�	{:���WV���eJǐ :[��+�k֘��Kæ�V�F�tVp����dHO�ӵ.�@d6+���G��g�粉�� �_�|Ȣ��w��$������؊#}�ll,�J��������]�>AX�`�t�/zp��J>��Αq���(V]���kmڌ�tQ�����7�yH�����q�b�~	mI)a�J���7��{RPoG��r�H��(�j�I�t\_Jn�R�hX��	^s�tV/�P�oZG�te�H�Q��ϔ�� �N�1��櫶��˕I�Zݣ�����_wh�S��k��Q:��=��)Ԛ�};?�聧�>L} 
�d܎���GA�=�f��<,t�q��
h֊��H8u�6��zd?�ZI[���7����y�����:6v(og
��)N�]�[%x��%n�eTJ
S�-�u=���eE�fѠ�-zP�΄����'�F8Y����Y3��Ѳ�����g>Y����P8�����[0w���o��f<W>��I���Ƽ��P��:��^�&}N�g�����[{?W�����"<C�$�W��S=�E�����k1��Sh��&y�B�k�yV�ժX#��b�����ďDB�%��'����=���~H:.��4����9>]}W�b���D�G�[S��@& �L��%���U�E�����_�D04p~��#*����s�
Kގ�yM��2{��L�l�����X�̈|��n$A��a[�>�E��F�)��]��&!�zkt�����
��8Bf�L�����K3��ک�9]��.+�5����-�����A��+��4��J�si�]�WuA�}��*�Nj��
�b�Q�]�Ꙋ��J�!���~��f�Y��a� ��@e��i+�R��O��eK�Pa-_6@�.r1&9��C�;K=CF�
��Wچ)N�k��1/��h�40#��*Ј���(o����+��:���D0j�^�t>G ��n	�%b���L�x?�Ж�E�=H��m���u��Q���c��'y���G>�J�epy��3�P�f��^�Oh���٤_*N��djs��3���7���d�y���Kn*�V��a�!�2��fS2��G�`V%��`�b�ō��-�/�nT<�EZ=��S)�LV�8����C?�6L�[��J�*$+
0천8^�����)՟�XtS��Ƙ����$ՙ�7v@RI5���[��UQ���Z>�k�|��'*\&�r��(\w�5�f��:��,����E:��,8EcF&�)@�����c��}'��m������N;�Z:t+�h}N� ���o���2,�S�!j��mc?(SZ���#P[@o%����2`8������ɂy��T��&��8F@��}����
J�s�7k�y�+}1��(���C�Q�w���KO�=�P]8>���[D�Q:��xZ�Emis.	a�'�Wjy+{�a�I7�3$U��s?w�xܢu}��T��V��od�m�9|ې?��;(+7�"K��8� �Rd���$㎋�_�3�l;(/�#�9Cr�&��������|J��p�!�)I}fl�Ia���WO=��X<�[���c��#�ݓ��Y�6V|�[b��C	���䭿_:��m��Q��c8�v9y�Q ��� ��P�Y+'�ޓ{�E烹���b,����j:�-�Y� ���������}������[��vZ�;~��D&�/�پf������سא�� -H���l֓�/����ŉ��� ݶHߕoإ6�Mb�ϱ�{�BL�s}� �*uXH���:�Z����$��al���ր�d�Y�\�_��a1��':��Qk[���V�\^`�Ol,�FH#{>~�>L�P���B:\������b�F�.Z	̰�H��[�~��4Z��Ψu� A������8\ag�겲&�2�Y�t�*�cZ\nɸ�1������;צ��\�?��\z�#{�[�K{�6�C(9e}~[Z�l�3w���XH����H����`!q@\��� 2�L�m���pL�z��g4D2-���n�9�iDt7��K%Yw��7�B�wl6������Av�-\K솬b�~Ĺ��x���1Zv��Y�86kZү�{Z�IǒS�m;K��>����R8�������ѳqEu�m�)n��Rq������] ��O�c7��[8B˶�r����!Q�����d��u����qEe� 1�4���Appq�w�.��$���\�p�s������w��KS��X�Njh��{G��Id�h�=\%m���� l/<g9=�ܝ�f-Co�B�(yGc|�S�c�O@�~���\�"jl�*��b6uܬz���*b4���Y7���t����>���:­W�P��Ոȡ�h{Ѧ��]�2� ��@?�}��&t�~C"$C�������p�#0��#�Fi��J݀�j���b�(�+�d�,��T�$��r�O�Ͷ�p��$�9KD$r]d�Ow��A�������fX8�L��\A�7������SpX2�?"\�ɲ�k�1�>G[G���;  i�=9oON߉ ��z2�"ׇ�����B��/m��ƫ�?r/���� {��1I���pې�����x�M�'p�:s�`6���.6��?��1{5��Q�ӾA�)-
��5}�ʶFj���^ٶŖ;�i*�U���g�U��-���l?寽��2@�ڽ5Q���T�ꡟ<�J���=�úq��Ѹ�W�X=�#Ċ�.�R�����1B��i(,���0����?���=�D�1!�~'.�w_{d!�+�r��v���=H���w%�(G�#j�f1=��Ωևߏ��۪�☗��ږ�l�t��i~98^R;�]�˽�h�}J�t5^C��r% q,V��F+FI|9|�1�9S�K�"�L���֖L�%�=#���򐑐ǌ��Rw�j���7��s�uD$ U��K�L['���m_��˳`�1��D��z?W͵���B	.��\^ሑ?�K�#ǭ]�'�\g9i� �@}Q�~v�H�l���G~8�������'�M�W�Y%�
sS<�z)��yE��I�+-0s���U�n�����j)����m��i���{���>���-*� z"�PO���5�]D�7"��Ȁ?𬖓�y�H�6݆���G_�F��Jyݺ�H'�H�����	��a�^f��:A����@�O&�{5ˆ��.����0W�XW����0Xv�e��	>H8���`F Ixe�E
�6�!��<�hh��<�ޢ_gn��ȯ��Y�����N<|N�Ԇ�!D)��"��Ϩ���5�iuS�5��u*̬��-4(�%R����9Lvc5-��NMe��������~�G>�PwJ�k4��ho����!$����G�1�i�Mz��n�_���`<�����	�J��!��2qtykuo<��_secqrXzV������Y�6y\�f"���I��
�'��f)�uL��*�Y{���2�H���)'�c�'�<�U$�>� w��Kf��E�A�t�2�A��>�i�kզP�g��ҹ%�Aݯ��٠�� �<� ����q��f�en����U�q�p�9�������j.��7����Y�/�m�ԑ�4��;�)c��Gr�sT��j�4ɦ~u�]ȑ�Q<ݖC���_k��i�mc *=,��SV~�Փ�
�K�������R)�J
�H���b�>�W�w�<t���*�S�:���kU�3��Y��_}�0���~/hl^�cu��BJ�^Fg�؇���%��� ,�?�w�V��Bo*�x8����f����P��!�0���RNx�]���y(��W�S�J!.�f`����l^�)��'n�X���0z�K��/z�10P��|.:�m�E��xw1�br����1S� ��ã�y�-X8t�:`�Yλ���:.x9�'�����ج��e;���;�����qRJO��SJ�\��h�p�R�]Ix$Fʇq������YzT�S�������)nr��BtiH˂�>O<-pX�P���y�ʍ
=��0�R���������T>���Cю�9�sqGOR�j�3��ZY�;��k�w�X۾�~�o�j�9n��o�O�HF��C���xJ�mܨ�\�S��%���=�V��@���i� S�O��/�a����N���X~i��(���bUR��yE��=[+�t�R$ �4�ȋ
1��%�W�N�'%��X(��� ��j����(�/\`x�\�ThD	#�	���pQ.�{�-o�U��}�)�<)��}�@����ʠ:�V��>�R��T�3�V{黁t��R!V� $ϡ:��b�/�����-z`ZۘUy��:�/|0		��?�9i}:���.�6g���g�H��H��J8	�3"�iO��|�L�F�OrM��H�%
q_/����IS�B��(�X����Q��������9�p(���Y1����V������	�O|�b�vH<�Yt�B)��w�,t�Ö��=�u��x�����xB��<�w�p?{��ȧ��)&W^��CݸGE\S��i<�O��E�\~��4�w���͊��G+�) G��AѢ�͊W^.�/�s��K�ב����$��jO��c��ښ��΋gP�B��&`�΀y�ㄚ]]9*���$�:�<BXwbU![�c��Fp��Ĵ�����od2�f:���*Y!�[���"c�fd��� �R����p�o�����-/��K'@tRƅY��Z�q:���f-�hx�>��k?,K����U���s�$��y��h�ph����6`�Gr ���uHW�3�xX��:�@g�J������V���GxÇ�u��78�� ��"|{��F�Q)H�SH����+�3؄��;�Z�Q��$~ZS^�D3P3���J="n�~��Y>�JC&B�[ך�-W�G���+�O(NF�����]G��]�`����U�?1��_�g����7	P�k��c�����U�$� ����Ŝ/���VT�G�
b	��삅�M�'��d:RF��ޒ݇*fi/�ҧ��&͙ �|�7[�ֺ��]I�'�:�0y>3C��i��X�)��VjN�xѢ�q��'����&��,���cJ����#H�� ��ZB�UY�|3���){ ��q��}�z׹]��:$�=	s�������:n�w�������VNB�6{�nT>���a�kh�M�1���e�n@9<��IdK��U^F7���$Kճ~���7q�'a@���U���k�rs�����c�߈��D��u.��;�9-`i�<3p(�@�g3��h�*��'	���5�=Z�(����u	��*Q*o<�I���d��a�yr��˟������t8�E�,���]�eՕ��+c2VҔ0`gɵ�kEpn�ce�T�]X�Op�NÆ҈�a-햙֢*D�Sa.�^��	����4�&2�+��0�e|~0t�G{Z�mg+�s��<��;���$y}"޴ �~5�P®M0��B,<+�,T�YE���֕�ɉo7�EK;�jڢq���N��)�/� ����,΢^8�/�H�|���Z�E���MD���4�A�F\`�4���� h��X��f.�e�uUg���Ȃ��<՘/�C02n'��)�V��'W�4�p@l}O��T_��e�w&����e�g���a�r�/���`1=��缺�7��]�xx�6?�3��5f�Ɍͣ�À���~V�hёz�B�t/��� W*�K���P���<n��կdy��i�w8�j2+ K�|���]�ڶ4�d|S���q{ih�K��h������̊�%������\�!,�^��A�������
�?��	��z���zS���E�����}��:s�_� ���P�qB�)�!����`���u�[S�r^����%#�޴�㟧��E�y-�O7"�eT�i��s��E��u����	ES�G~QoȤN����4��u�������=��:ߌņ�i,Q����\�2��B9&�͡�'�4��B�v+m��I��f�A_��,,+�J������^�o)�w��C~��=�D�r�3�D1�����YXs!دf��QF)1��9���j'�C�P$M��(��dl�y'�<C��S`ˬ����R��a��0�����L49��$^����JQ]$���p��4'��Nӿ7i
�sպ�� �U+�8e?��r%!��(c���4.֏zr8덢F��$��F���EAdj٪@)Ӻw�)*�/��y��oc? ֻ��г
r �K�.��u�����G��7�E"�5_�d~%L�̇�=!o'j�y�/�}��ߓAǒY�'h<���gz=m���;w��;(�l9K��&RS�3-��j��oy��a=�?{�&Ǎ����i�&����&3_�i�Eɮ`����10�Q�_�~� ��(x�V)�41b(���,�3� @MQƤFHQ_�?�j��+���϶-NB?��>��΃������Վ2Xe��h�����K9_�d��֗I�t�}���pV��f��߀�b��QxFgA4�aQ!�����o���Nud�[6T�����<a���.�S��tw�m΋�"J(�r�O�D�i`��{V���Qj'�����^$�B��Y��~Au:G_sX�gJ`\z�x���x�5�B����Ss6cC'�����9Й
ۑK��+�B]�3�UWZcE�>�x ya5�,�*K���jA4O�/gFW%ﯴc˩�^`��҅����i��pm��v�.1.t#�E+�ܣX4�ۋA��ϣݝW凙N��(�K�v�|�9��]y�m�;���Ok��f�n;���
��ϲ&��d���a���3�U�5eo��o��-{0�'����7���$A��oA�D����3�N����*����6�D��Cρ|�%k�Y�+�@ �t�{�p��*���sDB�t�С�R[bs����&N����jCm��[�� ���&v�r�c���vhQ��u<r��l�j�2M �2u��F AC���h�;���O���Ѐ������PW�ԁX.��9L(��4�G;�&�'&�26�B*���x�tx��W$��n����JQ��1��t9��{�vo6״MjT��D=���L$��1�� �2�@�Be�>���@�~u��EG�<�/��X��4,����pRJ7�Y%&��KU��KM3�`��	;���n3�?<��r��]�k9G�do�r�`�s����q��u�*[�⨽}a/��z`?���˭��7�ɩ�G�*���6WHǩ���^;b�� s��m�x|#����}������ؗ���X&N!ec���"*]��{5:��؂W�xǝ�ξ�j����P�Z�S�l�2h8�Y�\��XN�����g�cت�4��tw�Bc�nF�cc��~��F�� �l�N��G1m��L沌�;�(�H�8Q�������_"O%Bzf�֋ƿŎvo� A��)��u%1�����٣z�Kd�Q]���O�vx�3�$��l�N-�Ux�Ztro�l�������~��۬L�([�����C�+�NR�d�˨� OL���f� ��jT��L2� FA%��V��O����`��b�fV=�7����B5N��Or�]G�>؆t4�E��S�
��޶r�Tj����!&J�9h	��y���6�j���������N�Ԡ�`�Х���e;>�9�Gxi)$1*�g@S�U��q��N���x� �߼o|>Rfլ���V{"��Rhc�Ϋ;�%%H��P��G࠳��ø��Xђ� �0�<�Ƶ�<��"h�&�o����ՓI�cO~ܵ��-�5vH�0��9"aZY:��a#
�/���lK*���0u�c~a�I)zK:�K�T�]W��(�(��t+^%�"�pk����k���sVV@�v�rB��BT]���
�v�9:�\ظH*�\�P'	���W)}�LK=�y��{��v_�`,)1]�)�C4�n���R6m`��@{����}gjU{M��~���*[����᥎Q�bP1$&�|�Y~2�_8��C����V�М�y���A�loM0����Y_R�V������h��V	F�F �q|Č��{@abS0�Z�A�����n���H/ևd��]h���VpT9%*5��7���jW���Le2�Gz�ސ'iN���JkM;iP����ȶ�"�G�#�t��G;���p��B� S�tu��쯁�+�A�k�S�F
����r���Tho����f�Y5�?K�.昺9�xt8L��	�z�Y#�O�a<� 7�k\&$MK!����.�0�G���7���<��Z"#kb-}�A&wn7:����6{{�uwg&��.1��=S#F+{^G2�eD�Μ/Yp���y��VP�{vRz.Oz��O���+�.j�nVe� Y`�1 L?I[3�;���[�w�?R���&�7�ڎ�,�Xh�C^l^�8�fAW��^[�7e�h�t�%E/�A�qX�V��'�|X�}H�B����g� ˹J�:}6	����k�{XTF�� 0�K����V�Xi����/���h���I<��V�+<�����_Q��9̲��L��Fu��Y�Bʭ6�Ss1�+�Pʆ7RnhmT��%c��(6u�K(0�O�TF}�\ԕ�!���:�2�;���f�W�1~Ċ�	O��@�c[kW�{]������eR���s�!\��0Qi݈4�mp ۲P�e�9t���.������+	|��3���:������*J��{Xx������Xɀ^�:�����0�|Mj�ʎ2����"X<&��������_��b�&��؜���,Q�5��y^J���Vs ���T�l�mj�G�I0�@Pb�~6�,S���p�1��F��?�����p��ﶾ���_1�⽬ (L#�T3ʦ�m����:�@@�`D�F��\><Y��J����T���wۊ|������0ư�*]@�r^���k�Q`��3�+h޼k�`٪d�ο(ܺ졮�t��N����9S�xC�,�ԵR}G3��|�aj�{�q���G��a7.���n��S��`���j~�,�8���~Y}��L#�7���:އh�&탈l�]b|����r��X	wz��?�pbpV5��?�,W�7}��?�#͏��#��\��TV9Z��ܲtb�E�o�M!��������F#���
�+Rh��ag����ɿԓ 2Y?�"��0�i+�]��
��LgZx��JB���y]Y�����F�V��5H�9-�]2pG鯒�����p�%1���H�,U`���K���?U��x�ĭ"y�K]l�fr���b텸��%�ꑺ~�Iiޕ0�*�k�k1�udȮ�+̱�3�Αg��5��Y�_����e_Rz�L��"������_��;��:�p���e��v���DO������&6�%�Ir"�������ˈIog����Ԩ�Ye�t�Ft[��Q�#J7A����n������3H�2�O���\>�nB]U�U� K5�y�G�q��Z������)ddeG�����k��}�dK��'+N���,]�YXh�0M��h�~�3��w�>�����!�j�_f��^�
]:kK�{xaoZ(zZ!=g7�IQ�pE*�[b�'ҡli�Ӱ��8���8��J6�C�w=آ�u��_�w"�L>�l-,(��y-�5�	�/�~��L�hF9ܪ�c��|k�w�d��^������օ߰�cd/UgH5&����@Ԅ�~����nx�(����8+���1bؚ�I���?��5BI�{2n=�8�h��5�E9�:=���k�Gu�I"b
U�h��"��u|��ڃ�*���;���Z�E!�NMZ;�U��%o�ޣhb;�&"�ϼb-�jK`"f�NS�`��r� �n"w�ݽ4�/�M�|_z��36<�������G0�P���,����_���l�|ڬ�dC����� :��j�
qa��Cy��/�ǈ�LQP� b~���4�jF�4x8��@(������Jf���P�|
���oG|�8�N�h��̒���e/��[��*�ʽ~B�y���t̫V\��ֲ6M�*��z��1�=�~�_���y��C��`$?��@�a<޿xѴ��	��P���=4�L��h������>R��YS>�yxW�P�1��f$*�5s V��9_�5�